`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OBr+oOo5u/YbGu4kg8iLL6QTAfHxfOjuT/Agm44epiMT6kZ43/cKIuXcXcXJkRf4wRKl3tAmM4EU
99mgaSYqzw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tIlXr7xOahYPwMhLBLc5FESfV4r9QV/dweEKznRkLD7GhK+nKTeVQCyrdTaF1XYqT1KJDuMGt71f
ktSF14hLd25XbgHMlpswdY7KQl60mBuBoX4ytCyNplHo6tmIPPFIcVOfO3ok1HGNknpsIA6rFYpm
8KrN44HxAnxLnTsuZe4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kPJoKA2r7DtvguzHe7WXLXOtnqLCgPYE3Tq/wd+6MJokyhSTuAMVVZ+qJEXeqntSUAVRE8b5v0Cg
N5tt8bgopTtNRru6MpfHW0p5+xQVQKu9ozhkStvBeG7fTGM4yOH0g8qWcmPaDWp9q3UOq1zKlk9C
mmMEILZo+b/Ci9QfhAKgI1yVXy/6zJGT6CtLIBQ6Ap+XjzrOyuKQHbVqsUqYTwCS8Yi2zfR92rOg
u9fB0DuMf/qxdULDSrftiy3lZBHwPnDaKKq1dHcnidHuomTFu+oFOGxyWMsAEvHCm8zt5Ab/pjiX
3hAaIZz+/jXmZTqUGwV7s1pjDn4FeLhUBQq6yQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XYA5FRKSZXEo/HNS+eFDO9+jSq9u1KFpemZDrAj+mFynmVgY2Oh03xj+C73mfdrDnmUQiZAkjo9K
wx9w3TCU+kzYSYroRqs5XUJ9TXNhpWmYQEcGp4V+IUE4qDvm+/x5jJnYokLQCIZKSJym9+Ao/LdP
D0std7MtcqfXn1mQ+XI/RrSvS8zJLAKBT98bbkMqc9CdstWZvNi8e5srA5wM7ISlj0h4UWOh0JXp
8iRW5Vc5b4TLwz1+dTxaepg4wMOWR80LK4laRK3fGDgK+fHy6zIEHQZ8VssBs6c7r0PeHLwXWkwf
tBJ972k+/0avoRIbkj+yOVicvIep7SrfWiY9JQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
afdKXVTrNRiJjDy0d4UOOB/anPWdQGegcUW8IWaZ+RsLfCwDsqXaoH+aCjNn/WjgluZ7ntGpQHJs
o7pjzSdPTRZlmsoDwF6kDmdBX2zLQ31McqHD0vi+U/jLLcB3/2Q8Jm7vmh3b5UHrFd3ZtguYkgXC
6v13d0bNbxnYPHWexVE=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m8R+cYe+jSzJQtto8q1OFRYG5CaYdvyxwL+7mYJ1uF1crQMYLWNSQEz7SufvxVKL2euNPmaU5Var
opsHhzbMPih5qopKFRgu+ZRj6+UOUBNjkKkc0ueQXD/SiXZGSxvUX8ebOryMuWHDiSWMboNCSDHF
ME9XzMNjSfnqVhR3nGCF5O8rXq6YIy0mMmuyGlYHrYZatEy5fI7ZK5zkPpL0IYTIQvSNjyNEviVz
nh2dtiKLGr77UKkI6XKzWuqdtzyAj3kGbdtkFV2YdzMCih2UTnKk6xUGHhMe1dj0hfYpindg2gG0
0sa+AUKBR/tyR427giWUiVxTZJ96gEUyiexnCA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fmt6rTh3/uFvd2/y3pYZH3L3Dfydh57eEWeU2mWOX39BTs+vGsi/gYsZmHFA6ZSEYQUzJrlUM0Nt
aSqKglN0ukhlatfMU+I2oa72GfR31e4+jez9FsiaI3DnwAmdKJ1dQ0Kfqcy0qeSKTCYCpwpqjZui
vsLFmP/Jpecc9JdQ7Ii93a2ICPx+/BxHJh9IbJM0J9yUzEyElCeSPcCvTbjYUW2ylHUR/LKXtwm7
kxw+mB3fKuI9gi36aSLo/em/Qz8TckhsS4AiEBgVH0Vfnz20DQfCMsYT4I9/nwnqraOZETQstomH
Zr7GyMKxoQYZdRnQLJXImGIk2nWN1q/IcX62dQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W0q7R+UJ/sZjjIlIrcq4EZmmkrz3piz1O9Rn96Gbfdgl/3mdz+nwqJXGouk6Kx/esg4FrBEL135m
xFTLiGR6s3LoRF3QZ51rDmgp/HJwCI1HB9nu8TUdxJ/rThKuj0o3vHR6LUJhpXB+3SoNXbPfpLM0
g3dbiisxZL7/499rxG3tgj0GppDM8NgvPwnaP6+/OQjbwEA9Ji3qfED+fZ9ByO32vUnnXeCfqbZP
3ELzETUigGcqea3v1hgIonby8LzsMSdn2R0zobHWH+kG/UJ9GZtXHARewjJzizAqMDPZ9fYWuF49
wTJkKHhm3qZOs33x4ZRQruSpT3aIZ4bR+B10lg==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RMrZhPOyxeedufPZxYfEAv94x+xnbnwi9TXVGiAn6MHNOkuTiqD/0wDnuBYwaAtwmvtTqOiyZlKj
9RyXAPjxTlx3YJRUnibz6kzTyaOdRr3nsvbA17u5ULgKIs3BeJu/iAP2ViPFF+D9E9QOJpmmYbei
EeZc9cB81iouWnVqdTozJXgxyeZlzKPJWpMlgYcmm78tP4zsJEoDyZ/fxk6J9zdWVdOVX4SXJpp5
N/Rjf9utM3SmpkJJre2XKRXK6awAuLSQMAIVrXR5qw+UlEyvXLAXBpxswDICPKEfPmhcY13SeyD2
xEV5wGEux9qfAG3PNJC1yqP0Z+v6ywkNbh/V5Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64160)
`protect data_block
4RkUXFhJX6oLhAwDncQmuFdMjPVhY1Z0VT4MTbCDEKMWpk+xdbUBHD8k3ZbEna9gXmU+48/+6LKz
hpRYAjYFudBQa25MvmTincpiQrGbaFSBNy6Dl8EIAkn0V2qkhNHWBTTnxnzps+pdkz7ZW2bm0jJ5
0sqMnFQdyoN0HVjhOJqqVqK+nwrfuQiqpL3akq/Guv5aRKeD3Qxe0KHCInHGokchAv36Wid23QWU
M1mvuYKW775AerOZFVcZDqoebupiBvdUxvFosy5uLxt+5YgifvITgUCyhKwFJIKnUq8z3k90ARun
eyJv6u+TSzLnqhmjBlEpnhiZtFfFvSNlkmZLkg8P6HXi0Nst/uQyP7+7Z9Q2vtH4DHCpfA52jIIm
QglZndm7wBgbyRY3kGyVsHnLIlrozr+r3pIg/4OmfzWz2/w0BdMKm/qOMpOibJm09AA8A3cVebSK
XHgKJPMFaelEHlv16VKe0v36EIzXfJ2efEFoBSiNK0uFxatkZUAij6wwo+qC8YRbffEayW9te8Lr
6Z2xzdffRQYCXuFGDYyJN2d7OgIqAAULQgXRK1LWzAAEudSlhkp6HPfInB62+AZecWJNOGFWlL9+
ix2sFpiDv3rU4De8wCwTBE9caRier+TGrgvU+2wdKqAld5L6b6ZH164wi9Mw4heEXl3rKG49inHb
dmtr68JUiklTVb6ssyh2u5/baBBtl8AFzehaq8NCaIhR4uyolNI79+9lXMX8K5l230jhIy9QJvDv
iUIJ6I/MEgPvsA0GlRKs8XycUZyEOvzrrluQx2le9fGDemMLSMFGYuz2/1yv6zRI+CGuguH/lBkG
yxqUVPSD2u7Er6LVDbuLm6z9z0BqxvDG2MacrZV4d8bnEDkhk73qBprkC7RljwGDCfPXx0cyJNIJ
IbZTHkRmQvSZztvvsXp9sq6lU1/IsBinlSGpfZbINjhA76A3I4EgvYBWBQAEqw3QZ+Y8EGTerTaJ
OSCkWzAzuKV3ceAsoXnCQQcHWk1+5V7VpBHPHMHxSpO9j2iRzj/FIw5dRQI44i5sLVTyVa7C9fwi
kj7zB3oBflomVZB/TCTnnT9NMYyt15mUosH9K8bcK057tznN4WhVWwcVHjn1u41NqkFtnisO5ALI
CTZLyPneMr8YNFht4LRgFAHJoe4O8mGuUUPBldOt8Y0uW4owpfytTToIrnDpkbjSjGlphoPMkX5T
7labCu2GKc1pbf2EkDScEAFvzmg05JU6Q/XyRtiiXj8R5ha1VIZkZ4EBtHhMewHdfKM8MKOqFXKE
gIOeZLY0h7Ko5bVod445FDEIAQiQLSbDJ+hRcjYadKrmv9tUnP1NN9HpDj0tHKoyJ9LGaIrr5Siv
fOAfa6cN5c6jv9ukTacXxP7mwp5ubzRwpXile74ZuKzPq2rjV+yjF5YdD5Xyfjvm5gVXXcxQHf/F
C5zSxeGZdz1NIdwSN9jzD6VeGq5AdCykDBCAFD9xEVYhILw5W9FNJCLJzA7MifUH9otgw6uyMYwl
qtGxKW9Op9RHlrMe7kQjSLYZqkk7wRJDiiN1rlsNnTvqisByJlz+jlUlTngsWXVk/ibi4AylL6op
A4Uqdlpg9bzPvWDjgUxMGU+O3gJoN47v65MCRM/XiHRQd99TMTroqrh4eZ3yj0pAPPqL+7pSmLtT
mssvQhDSBT+RaNi1dq9HA3faKpHEY9bfcvN/1Vx5ATrubftiV96N3FUqtHjsVdbwAvs10mpN1O0d
R2NNcUFI3VvAMQobzEoOVHFJhPrUIoqHgXviRN2Mrfk6hR6jdeDD+VDdbTp0VkvxQn50R2jFME0r
2B/kL8zyQhIRUi3BFOAMrmofsYCAh+H4PYrsmjRlejOy9fX33wMDKLonGQhiQd7D5fwfzm8WVD2c
DH/vOHkEshjgcznci4sowyWt2WLXNMAb4TBoWbkzvpIr24ORVtHWdK+9sqHGhUwYAYt1voavdboR
kNEi7ahuRJVgC491avRFXgNjAXE8U0rjfoSCC9l6IKEEVtec5V1pfhvULDgl4u7cpYtGFcPcSF+d
6NGfV+3PM5Mig08dTVcub/yN9WhreEs+h1HBGrauNHh1HuOc4XuBrLJU4D7szPknqJp+iiO5mL8K
S5vlmIihfKw6YrBKCR5OlyEpj2No+Wee+KJRvsyyhTp3u1FSD/bG9bIXr9mDV9NAeKOiYXPGTa9u
gKvf7WrDWEzgsOeBo14vuDEnMOYAejROWD+YCfTuNIcvGYduullAuwLR7wPIs8hNJ08L4aFWfE9e
9N8Z2Na93lNv2V+PVNIZDpkH13vJwXmUJcxx0CL/6H1AXfH4TCyq4zGgosovqJARa5/LXk5gmOf7
AS7IEsQ3lyhLAcNlHl5B+XrA1FkrBM3Km2gDXwZgm/q6agbY4gC9T1scalBzaD9xsGeZQ5rAo2VM
Nq6sR0AH6eM3GpCpDo7xGj8NSD0Sfp0rupkbcx+txHOpdPDzR5TLsYMTeWAdH4s2S/JAEv4PRGqK
P+Kz7v9nPG+/FmDIPAf+0zGVdrRUzrldmdZGcFbsv8j6C8hnYIBsuNDul+O9TycFv0FAJPk42bW0
JD0IfNKcwJ0wvBWTZ/8pbkgNt7UZeUWC6bmyZblW2rYk+PsV8sJU6x7FhRJGixOx2kMc+k1dRK5y
bTAOgv1xWDGQXXBtVkCCaGpy71n8uxOo3aRjYMsAulz/5WlC/VvWohpUHiXRuxcfzSktw445s4TC
f8kK4fsWC3uOe4Op9MK+6UUf8VjztnJCQmnvl4YAthXLvIfh69rjxTMdWdJjSPzEVczo7AERPSSI
6kEzaX8Uj8X9KeuYhwGHz00nFU5hOyWH9AAr8PfkvyDC0T65zmg11VJ1oPf9hHs6/a64dTDKTtd2
yb45hLhbngpi9uAhLzz9qRDs84zng1jPwBgdsMXRLmdXD2Bv8OW24vBHgAev0UmVad5QGgMP0ojR
UJuy0n5tJVpMWaXKx1sgK9H7JNtDmhpDM6xZrgXopwF8JEtDNv7lMZtCCs4OKi9L2GzAPoX39eCh
m3SoXF2MQ2q/aF+hWTpV79FLR0oe4c4hsXEsHBYlm+qbuWMjvFzuLlTYZChhorEy0Vr2BWY+5KJ0
G2O7lRdZeLuROkHJzam7H+SDbY5/ykaOW9OcuU97trbtyeePdGwn20YDczB4Oz2J3xo23jl+BF8w
Bk3RDRU9VDpPhahetbQd0N9OM/4KIpZ9uGg7CaoVIF+i4MM2Wky7HKAD19ST5u/9aGliexgumfmY
R1WWdSe1+E5SLj8iJID9EJLqS+YZBVMzHPLAcWZ+wO4mdDXKeyzbGkVazvUHW+I6L0jA/mezFMVP
4janB+ZyemTsfmNQGvId1SAb9kJwJSQrdvlCt0KknlR9I1o0sv8KcFeUl5qNKaEUqFHkGNZCc/2x
+RC3EhKf+JBWF57QP3Fm66uhUu9zU0YXcrCor+NGu2xCydsifnLL6IOSi7c3A43rCA/OjJpzsREr
+GiB0qlM9dCTfd5J3m65CHpH/dR0uPnQcd+YT0C25I9p+2IpAFlIcYWvyhg1pjnHEpD+j/hnZ5m7
9z3pIWfZPFS2gFF6Gm9bctq8PTcHjfKywv8BQFuB9uNADtGAXRl2LmDLsYtrWDqwiN772ikJ9zQi
1WxYLq7EfypvdP8y6UOuRP/VOptGV+pqX5gwNt2N8qR9yPpRuiW+MaJn4bW7Q/VhH4OH9KMSteXH
3fhHgtBX7txNVUuPebap2eA+jb7BCPiDV8I0854Q2Rvj6wIUMvRpXGG57tmfrVfovoy+a0yuaEhZ
GtagErp84MI8Fg1ep3xVvBC13SetNcqjrP9x2ySikC26u+Rc6VcKO1VXEeLUNOQNKDxc3ZwXWeY4
0M/RlBo8fmJ0zcT2fquRg4tDDnoKijEgnpbo700U3soNinA3Ta0eOtalrg74OrNoPkdNX12ZReiB
YUpKNdE7m5gcfQot/vT4HwE0q1SQEj0AQb27nYm86d2ODih6HAWZuU40pt29RLW2OOY6wfaopANl
9rSpZ2JAzLL3STn9h8D6yrBlNOvHjioQmd5aBBKAX4loa4qONmozK8eQgN+NjCdt5UsT2h01yACk
R2JgUPR+3t2pRdmJe2ItHfW1fn1QcGW2iG+Iml9xwgmjrhbKeuMeLp57nFPtWEgNqRKsV3mdfELs
UBsktqprSQHDWmxohnUhXXCXd0KMCv2mKn7mXmBSjmmrInnVLnjyTnRgDR2JuKS55AqE2tHsSDdj
5aFiAJb3QfWcfV064/r4t2kCjinpbPnEtJGn+1s6KYtjfT7GW4BvGdJP2rSgUjVEJVFpvcb8Jf0r
j1N3F0GPMg9szheh9fXdf5f/muQ1yE1WN8D5akle1aqjqDDAk0pcwT8EFtuyol2VWCIWBIsuI3kB
1V/m4gi7xfUBCV6CCaajOyni7pPBl/zuXb+K53ku274GBiDCQWr4+GguxZ0UGdMhBKBURHHMX1+Y
jpRaHaMA1k0vM7TEHZBPA1wptjtuEd53yKENMotoCNdzNqdXEIloApUKk2Mj65vw3CmDH7Jsdprb
XO1F8rS3LAlvi0xf0FFNpw9bqg0/v4U5fN/lOwEgPQ01ENtO/KMvE0EFoDqrktNABFjXF0y8iE5f
IS0SdPebDc5O758TnA3hap0jx8zZ4cZ4NoxrCqNrrrkCPsocGc+NhLXwZBKzLMPkaY+t7q2huotl
Lc5DH1lQ14wmb13CUCKO7Arh092IrJzuhBs5TkGlWHIaaDct5uE1xZ/fBzu1+bULuCs4DXnKieaD
QLlle0DjpExcs/vuunQHszLanajO/UIbCVLijYmXf1BIya7JNeaA3Ztg9mi3H0GYbP9olgMtoFll
G6LuyVmmk4fQApF7bnREtB9AI9jzduDysLJUn6tQ28IXXHfiv6WvhIaKRSH0IvWQQE14oTQLC+nf
poX7pYdGNKxYwCvdchSUDsJi5Ff2LOnd25BGnYCtCDCEK14NzfqmP+Xn3D8i++2I5Hka3CMy2X/L
dWQC0krwgHhYj/qbdovWHC/pvk9kwFxm8AMaMhZ/ub1t1AYN0yNin5c/S9hRBYlDvytqX6JSp7/m
m2pDx8Q2JX0JSIaphiA20NWSz9GL3IVt6zJ+RvsUIqX573LxMDzSPltHF68LUseWdCccZ7xBSc8m
7EDdz2hQwEKc2O3Sz/1bS1a+r/h8SY7OF/OsgulDGK1NHh6cA13C/FdRgeT1On4iRi8SLpcTky5m
wNs69sM1n9HvbVAsrXhCJEWvq0q9LKT/3FBV4X4U/cZvU0oDQEsfbgzlaZUwtevzSGoKtRJ/vAcG
gurAlCKvuXAt13L+0Yi7LOojhNTXWeZ5CAQ5+Sic1eFccl4lBmOmEFaXUMvUsf8wO/R0GGn+4NMN
sALsMaT1iIihEXCCVnPEWJpi3uTyttTAn8QLAVbrX3D2mq9qTE1HCZJ+K9+TOmoWC79fsl+V1jZ8
l37NiqmT3/XUvCMVZj+w9k59dvicXDKX/fJcgWkj0oxpdyZo/hTEBDjvvwYmSo1XHWmCzpw2JgfK
pX0dk1JJHk19o7P5SwP4v04HChCfwChqMnkQaUZ4vLEKZ7Q+MvMHhy0IFB4MQDaAg4ybd0H8NB/o
s0gQRjr4mGZkFpOOfZkIxV+Ty/9gGBhPjamAX4vLRuwwPyQXaMjfqmaLGQE7wCvHLhPR1C6nlS2m
UrjUNumSban2ceJJtsVzvOi1RZQgGq3c8y3S7bssoMkckBz7FXQcdTP+jnX6/8SWTS1qQIQS7yll
fYrBR6poexYDBKuivalCa4XaggMHC5KEHPdE33Akzth2HBRnFX9aVix+roQQy1/UKikJuYWG5jEB
pe8F9UoF3h4jgaF5BxfUkGePPc0pNcpafPtqrxzgF4NNk1WNutmpfuVQzDrgDItmf2ncx1JLfQBk
BPqSWu9vPoNodGFx4mE6l8DJYroJ7mJ8z1xT5xW9SWqoCBCzELNSnwOGZbsuNZGfWIQ4NesHBQX+
I8qsNkGihCPGd4qJUPzhFmRKg/2KxmXHqKY+ARTp/9A1/MIdqMhf4FV+LkUlc/pCsjFHL+KLd0Q9
6bLpvX91qfptGsIn2ddhjHDlwtcyfg7HwtoVLOr4x7o8oforVHnoZYYefYqx6GwJ/sfR72Yg5PdG
UIul4ahLvgMT7QeVv5PP0DsXVn0YQWn8ows3IPJcZyAMD3QXcdAHa71JRfc8o097rwF8mFDb7gFj
pgUw+WX02JMAM15OpNezXb0kR3vVcz3E0odB1C/MSosZNhWqgkcl7hoj37ggCDZIIT6LbuXA0myM
4M+PQpT4xxVQWYI0s+iBRQlF0IIIzLqDgY5pxq2DYi5MghaPDodrqL8PcEoplgDnI/Lz9gC/dtFL
dyEpK1EFdArl2k4jWEwHNL3RjOD82JGHbk5nFwVBekTevlfi1TZifhukGmn+LioHwzRD+WEoJG3/
+G3pf1pVnZC2Pfbst67sdOe8KrRVzwoOQgyH5/le4EQWV2LwoZPxjIbFHrpcQtBU88xnPYFDs980
1Yp0hf1lDLCXKduD2RXWKfadu2/HIiH2GA8PH/F+KkW70wPBswvg3tQJvhXumU3lEtUluAgUdf+W
Vrau5WPTFoLR3Xsu7EV9R5gTXhDs759UtFhFeSvskzShG/fHspfDLl9acDb5LV/xHamtWKAdHZFi
0+HYJaCxprOxpEN7m6jGbdjFQm8tQdYLgJ0NKvIgekhwKFJDkdUzM9zgJiCt6c0MePLLFXCPi7cP
OnOP5dtuWwVxh43QKTytxY+hbt2HvfQMflEc2d34BmkuIwSWrMqXk4IScCzmAtuoickkwUjHg32S
f6wLGnuOXY0BjsUtQbnnpyB1HJGHlrjY0Afst5AbNsdAuBm3aHPLMYt94bq9SL+SbNtnwdIUJgtX
cPZSw4dXvLWr8fzvWIvq7Ers1wuoTnqWWGnZorZe6qXxduSUIOcVgMyKHT3RwuC4ekiJq/lFkOZ7
smQ4EGW9UCetAQLtp9ipiAsG0t4EgwTQ8cgJsJOp3MEmpeY7ZoMYciKwHPCsoqc/+uCvQZ/3LxHR
8UrInRX8+GVD8+YdykUuzllcUGrb5LzxOFWhwXH6WrWneL03dVzFx76eLiOhXLgZ1BXBXtrUIh/y
fHXB3l12queF5WLqIOImYIvo58uzNhMcnnFZvr3ckn3ph+LMkaRnjIIJkXJLW2+rff36tC55dXT7
XivRCXvHnTgILP+HI4c3ENCQYRe3Nl+/vLg6qNsYsI0p3Bp6W7MigNFuXMWR3tVnSbOjY7TtfUoW
vhvzUcVcGCCWaSvZpLnGTvJXwGT+/QJXBuF/MkjSNyKsFvi3eCkCvLRV1VFe52zuUMnCFX6PwxBx
E4kRjZYoUb/U2S9llawLLmdrXlcPZuG9vTmVOOrZFgzZOKvm682AflzSr4SRkgUUkjDQgPJRdOLW
qYvL+mfJuT2K/ekRyYoDQZ7cdFQXFCEfNUQxgq9HZ2XasL/hG51C4hCMo9KOsuX6YLUEiVlNguLG
imDis3u0eVGrCOfnUFdb3RT47fmaWgyDPbWAEnf8NXig8nui4Onos6eP+4O2OeW8lUIbKPB7kmsz
iJrcdl2xsAbH7DWWFrEVwKB6SgibJ7Cn32AWruqICV1B8KAXDOndXJRPH9/9XmwUm+HXp0XpqBCu
Pfkg9TW2Ja/jQIRi1WZXb706BcQIODU9gmEXKFVVR+t7Ej9FNEj+8+sj1u80u9CwMzvFJ7T+NIiF
1CUbwyE/0NbD2Jc/uPCZZ5+jPcCpapJnrfXhzVbrdtU0auR5ztciAU6GPNJnBf256I/gU5I51WIl
DFAVvIbHF2TFmiMrTQRWbzuefZPIkaynrzwoZylXmIQVMT6QNg5OQBuP+og0TKgpZZ5uYwyhgi4X
O8EXvAM+0zBBkhcB2y/NXZxCjGDiU6DEzF75MSi6o+DJiGfCkIwKiIFg5uKTMQqWfi09KdH3S41u
KvMznm+fQbxfVKELSKTO5gynay35wDz4sQlSRMqABQVWVzcbq+xt1OPx6dkXoUIhdDDO0inKZ8J8
pXft9ThyyAuWQM95VCEc5SOvN0LWi3KUqpXHvCV29EYpyKzCqntoVWAujTqkQ9kEBqXOB6ikw+v2
y9olM0BTkgwU6YKcsBZPnGsaHY1pWZFrYi/PHYh3n0wsnvavBfFUpNSPzDFIk46zbV3ZCHwJJToP
hP8j+iUEBKW/AvuiHpkVvnPRVL9P1EOxxrQwRnzw6h0BOC5s4jQq/3SyRz+8DwfQCrDv8YSDXGF3
HEBMAuxAUgaiVefYojxO1feqzc4yRf9dgAj/rt3GU94tg8/IVhomHKI/3K4LhX3PfA5VdIyXi/+E
d6wo9ygwy2RSlw4YlgFHyKjD8TIYRoNhNiOl69C9F4u8APhETXKwQ58Z2Dq8ybVagKsda7NtDEMt
tq7tamJTOfHIDgGRLeSit+XQo+aeHWUCwuQm6w86tAghJmRz6Ixaf2clLGb/FRJ3JrOdJmWLMVka
XpCvDX4+myRW9NEakL7bCcMGzBx7RPaFPf5fyXinxQ57bbMkEJJBggCFWvjnbyTlW5Q1b0xwaq+Z
dqassJFm1E9wM43izZI55zbrAyQe7bRJa3/8YyK/WdgWJrwY7SNlHkmDuZ2kJ5hXB1nhIbOkMzsK
1zyh6Q/9PTbSrkXQvY0VRWDTfo2QiJ2ckf1uYot1zvVJdSZQDFaJR9l91qJZ08jt41syKo1twp0J
XPmu4uyzrtpVv2kkw4UfKZAMwax0R7TNs6Hvcw3AkLI+hhGrXSZGpw+aj2v3PjphiN4O45MSYiKp
D2I/+2OIXDKlp3qwloCUxGtPeajer3wT11xzr1UNcmAoGmR9XiRmjdxeJrvDoFMmtPqT/MhqMlPx
SRMxIW+sLv8YlzBygSr3Ro8JQapCVuZ+2z+rEt9zVFNCxSVn39ZD7QWovkvIi2eZ7yO++IeOJcnz
M5i02Ge4QavUMKPzhw/dxVMamlfSqsnSIXf8jALLeeFe0yzfjLvDB/y995p+agC1DQKY7vx2w5r7
PLKwodXaPPylpdCgPGZlqC9SlD4Ml9fMH2Q076/akMpGPTD+wfW+pz0R9mzOXuX9+cEry7pDVvon
IwtgErk+RR1M0ClkJEcBoMZoDGCr0xqzy86wUqsYmYAG+8kFs3l9MpxXwBXGWxGP07G5otWTQAQJ
4LhVONCeJOagy+1a7t1flULA3qGhKRb26JPQvM5Vq8Aw39jpDayh8S4VgOXW0Zhi91xiupY0J3Az
R4exsn6+p/ygpRS/JZIHhCIQRimWkWqUxIHgOj9aO3cK34SQyo3o2dWB+QGY8z+AaDi5xXyQOIkW
HiZsq4SVFZlZX8vpoQm4S6QD/aabfKcpm/fq5PhZwvgksYH2Ze5QfUZmjElB4ISW900096LoPCFv
CopUimSBMe4sLYVr9rApqJT/2vMCTpF2+wAMvOJ8a/iZ+skC9p2qJpWoTsK6ihcN11qG1R7NMcuC
ur8sObtSp+wCjlEvJmRhE5HpOEDAdx6y7qRg/799kMB8VDZB03iciEgEmgxUtGnE4UaMLZ+6bT39
6sBiw+U+BAAJg6vIDsT08nTsHmMyk+nDkSnp/lHFr4YtzC2G6B0BmWsEBatSw9hCgHQMYdw6aq7q
C7FnlEiTLU0ffK0PiD7VWm168Px7zGPAG4yd2iH/1/t7j12FW6TrsNfcS1ZfkL9zjLGbHYwDf7R2
ZPyAwtvyBCVM0O+ry998SBpHUTpIN3g3wEvo8dWkY3nakjwgDmGIeCkWVCGK4txgGM9RWzkblOau
PyIx840i+T+uf8fbkdx1uT7KnHtrTKGUFcuWhVnkQcudXtumvNMQz1qBx3shRG+9EA4yiPKKwhid
C1OXbm5PDkDFnpr1ktzUA5p2Lnmi47NzyYWl35MWr3yrdIItDuTTcd+z/Evzm4H8OLb6j5T7cYtB
MsSps2vgYEIHhg7NUouG2j3dbqfpM3Ev2fNvdw4Rrn13kmVabGTe/mmYwaK1cowwgOXc8jC3DXrZ
H8YCwH0QXr9R9EwrgGZWD9fsZ+iEqIUiRX8i4N8bXlpwo1jK4BQMYDnuJE4/QW+vFlqf08f7GNTW
TNY3qni1h/Kw8XYPeG9TLRMMP/FqcIAhLr6BhobmsFts8cc3S28NUMXcl2iQHRfOrbYS4ueVBSDA
UmcdwtaLhEMKB9B9fVYfgX+NIYs7V7ueuYfVJUBQX38sXXUtmpuHtCkpHnQ6LPzuK+hUFaCybO7o
ogGSOp/++lsnt+UWQRACMJNp5Nmh02MLZ/Sv6ipFV+RpDicd0lhfkoAAzKuo5iblz5V0ISj7rvQC
2hJfX0Fu0gflMesZfRC7Va3OCp/hZvDKKZfZtFQKuaOohcFYclKD++PFYG7BU74937aPj954Smsi
Z7aCJ9/cuFX0I2QY26e456pC9Tlv/cxn+Bkce5iKvCSl9HR8JOR0CzJ0bYNtFcqDdEDbMhSV16mr
/kQkziH7DVmGuw6GumtMeuEWZt2X2OE3XsEoqYeHDWmIjztaa5RIVWN2teXDlZOjQ6Wirfnow0qK
eRvJ0QGb7ze3siNf3hv+BsPRl/2vqNhYCdYno7fTh38IziI5ADUfUHGq7h4k/RR6MS96ipT6c87z
4gz46fTij9BxMxMUZB6qil54j8l8lF9v+ltfLBlTbS4nEOB0BEcMOaPLedVZulIVXq7IJs1M5L0T
qqOmMGt2/uQxMqG3n/zbH/01I79ifDt5eLtywMGRaoiZHH1cYp3i+HTWs2D0kWSmGobzAUpDlet/
PEetzvU7TmhHCY+m0MN8NeE0IJpYgWS+WWLjE1iiHC7T/ieE6Xk0P2u1vOBSHTsNUQjJycKot0Cn
kiiulXDHBejxeZRro0hnYwxtD+3aw0SwlBBxXSbY1MFzESVKYXiEmd2T4vV+J+h06gJgzKFmTLYj
jqM9FeY68OYNdMjgotYiRs3rGY/+pO3Ge5OZH7kN4CJX1akELiOTIdNmS1GSK0XxK5eAGEwp3pVY
wBrjBLfoUp77nXhvtCz2rUIx1khOb/9yGIy4rTyKE1CMjjr4SPilzda4MnDy4ak5LepST7TJ9aKh
86C4KHFkkfQkwHxEKRstnbUE/Ap1Fx+i84AUXwJAAEhrwhB2ZsukUIjwTKdF7HAipAmjeayFQsrP
ePyaGGri8dR7W5RuwQD4rctfodqJHHrLF5PWASnVKgGr3AMnFzFdQjN8iZ+yoqI1xBgLOjB0dYi1
diSEWrFA6UiZySaCvOiiDZ8xeNhCl3pIDnlixe9WjUSTJd7qeRhNFXYy+103ste94oT1Gyv+Eey8
ZwjhAMPEbW69IdRqoC9MdyP52+M14co+eE+c0navkNiZlxHiIAH283zauIO9GMKZuVvFDGMzUtbD
WDOKaUIrzxhG/3fEGFZ2FhTxXPHqnbx4AO8IfjlrgMMIIDg2zemvTCo8HtN2zBK5Bpv6S3/zWPro
/ZtvoumjQTOOtajnwteC6RnT1H92bMjMLltJH4KpAJy6+1hTEbYmviAMlauAl0Dtf+zyODYcGqVR
6s4n6UaJiR30nUFipWC9PBLOH0z2jqU52j1/fREPhT7Xb8kSYUipn6dyuDJmGmKlsQmARm1Mk9oV
m0+Jwog15l5ayNrWkDLTlVBswoQYz7xw0+l17jE3I3AM5NNXmYuZC3y4IVLBW0Ctm21MMNM6MruJ
mm/7Dn87P3XRV9QHoAqB81sQQbPGk5OW77b3MChdL/rP3d+c+zWji1OC7Oh8Q4pU33sbpSnWriWV
hggxaIXvlLTIMGNvX1tkctBWuI2BtY5465rMvbOIwAL484sXHphBU1KI7OxEdI8Kubg1LfMyyUnN
RaJwwxGI9/y9BP5gF9ZokrvNpTCFJPOVi8W5NJRUm3C3seUJN/Y0ZOXNoQgUAfJeqab8U44l49oM
x2Lb+vH1PbJUkZIOqw6UBZa4sv3rqIQjwmFeU/8i3jztYLUpYHTQ4N4NxLEWESAVYjXc2BbU5ZVF
O/uXTnO2RJCFFm7QCoSWQUUOina7SbYATDoXv9UCf4dwq7cUbohDvbfjT2iX9c9PSdgQ5HAzjgw4
ZAVAplmo3bzVO0FHnuSJdKPlmnEH0QpmfCXFrWxCZ2bWwvJk1gjpUjC63s1mLNmHyTdgISi5fnAD
r0b2Zk/hqX8ZhBeobkFvwhYKpDiPgkr7NVGWHnJ0j7qOd8X+d0cYrRSuQOD2EaYTw/sFPSh5rVue
cdCXLpOdqhaiSY+OjmwmhxOHtgiLVrNHbpuz68gLGsUK+DMk73FXL2V/HU1TyebyJXloRnuoNqeI
77fC3PU2Xp00e1QwgjZmaLrrdOe84dNthRKKw8ZjNlfmzch2KWXL19aKIyqmaUfqMh1Rg1V3xVQO
Jlu+CQgB0U2oEK3EDlml+eda3eeJgUPt0fY5qKII5hSM2l2sDAKDphpUIK30274keatz+Te8gElw
+VOhMFQZEhWe7VGI3HEdeOqhKnlpvaVEbxNzRCA5jofuJ5qTmdF/4jOsGOekntbhe6zdwrPT+1RJ
vtNXz9ambVoqmIvm+/nzKYJL3uBLAkZYAoc/lx890YBCcic8o2Bn4BDiw4TTOGrSUHAv/0EVDo8B
x7qsNUppOO35zRhm9WV++Yc7Q07oION6paQ3z8wBNjqBFFR1SV5zyxa+Xs2FI02PrFLsorQUHbrM
cXR3+eSsDA5uZzSvbT+vFUwp0jeLsuDUsDm0ElTnI2yB5Nw56umYNaUcCybJq7OXJazCdPJjbRYV
a2CRAH7Xj7JsETFCowjvdgKtTprZygNqwvL7mRFrXsc6Td7gmzYKiliR40GPSTvHnsUbcEzwEaHj
u1N6Y0MwE83NAaPAKNA2BGF2tblIqJBBRzLDmiJLhL9lYtQ5K0oLccUHJmEE39fOFKJzMZbL6OMk
9Dy2y6OQD3sGcxJXyUJe6poQ2EpD2hbifB7JytZ4TYHPCUG7GxbRjvBfODrCqyR/kihULqpVAegF
HD9CUdsKFUkEDbh5QC8O3XuEmlnW0N2oZNAf3mEY3mql/degJK7bB5PYcMU50m6lqPK+buGIZgtA
6BpVIrvrpOaTQFXGMwa0bnYiK2iMXnpEdJz2ysfZpchPMrXyFve7SXfcnfNF0sfgQYmNc83wBLVV
4iOW3g1Wuaw263Q3/oBKQ4RtCF64nqKQ2JbgzVLjWmTQDWyM5dukBWrZsj6SVRMfkFKYaIxvUYYj
8q/F0UP4SlZ537lZ6cAiT0D+QBw9h0u2+UGI6nqA2IKJtpmP/5sthd2gAuZxouUtQs08g1WipXvj
oSJQLvtKMtQCOpAg3jC8Fmxkj1rgcjf0PE9fJij4o90xIjGAvmu8OIM8m/6hFfo0iP5JrjMFg58I
hGzC6zYAtyxEEBxqWPYVzqvjoZt59cp5NTqQau9W1Mv3kr3L4SLng9aO0qk84sWbfbmAgLsGjk/J
saGDaA0hoFFEed01PfIul3wJSXqvKrJV0WXh03U99DoYkzLvhyUe8+kKG+zgOWIszzWK9/rlLrgk
7MjkXVtbHwmzcfWSuC9coWQWDOOkPlRyouq9U/1BxKyN/0Svrlqn3H8rLOuJvjLvl/2fH64XHCfs
5EAK/pvv3Hi1tKZL6ESWDplZGF0r6BYi5MGjq6j1f0Zt0UZToXeyDMiEeXr1gHL7pn4ETEbOiytM
BiB6ipMCd4wGUF+Lf9TPDNBWXYyG+T0T6zNr4ifIE7+Wqr8WCP1cuSiQsl6mj0l38Rsi/tVPzaq+
PoPFCuoSJwbRcuCzCTtYpvrxQdLN2785EgE2qzcrjarxY6pQI/95uURnypAwjyFClJoG/NSKxn4H
1pijYV6YtD9svnEGDOKYgTdtIq54YC0ro0kj2CFjj/j7hIzllqsmdTP70LT2DFuFnYOXzgB5nzK8
QNM/sZRjtnAElzLNz3V6eEW2CzxrAYaFsh/g4wltL9yMfcU6WyBGz3tqMZ0vaowSj7UqAODPrjRX
K49jE/SZnJS5LGxVpsWxyIhcfvcg4pGyK3Og2LVmb65olA1s4LhzW1BeViBCCwSyMr6XBTksgTon
51nACkArph+ZFoUQgePxxWRPs/hHSW3BUSQq43/RS+aGhMZK+5e002/4TkPuHzNAivZ2VQ99mkaB
FpZ3K1V4qLPczpo5pxJZPPSuWUcwOVFnk30cvMlfLhTDdDZHseV7E7m0oxMbXfO0p7eUKejcwVYz
UDO9f2TQ3jberzjRLUoh5hLAJontRTSoSR35PpYUYVnc2XYmwSGisr2Rh+vAo9nG8RzG16pK0ytt
JODsZ1lOsFpwzjYh2sx3IpcwcaNDeaQfpdGeqVM8xtsaw4sOLzD2RREXpmyNwxJLIK0t/En/vIRS
20SCFqA2zbdLOnS4kAzCkT4j8SryEldXhFe8mvgl9+2JdNvdm4qTiCl7rgKbzNQgNJmRmckFAANW
fDMSRnH0Oj8kDqtwdHXHYQ715HuawgNTWjpy+ox5hqWUiG41IUHcU8jKUdLAcbfKDG3Vxu7PzlZ8
p0TfKcFfO6NyqSLzqfmv4XafG748OPFx3+E2LNdCrthMMepqGbsnM2pOoWpzcZqT2Y0zQoQ+ktdX
XCc+4FsWfshJ0q9tfCtrWvxbibEkvAvW9eQQE/tVxwvhZfiNPmaPp+Xj+bwerZ6klB63cJuKdKTX
zwEUL1fsyRddrYPGHr7x+A0raZzs7S3WH9VQ4NGULrUpl+ha6XdCHYmSFxAl8A/SVS18QGe5Qics
MOg/WUGicuxn1xXJ9FcAGRQs6OlovdtJMsWzpguqDPEdFBIvhhw2pSBSNTQ8uJZdIhh1T8XHEUAU
2Jy9ounvcpqQg9Z0Dqx2eWHAMNs8FkZcoDywNltWMdlW3O+uFS6r0J8sXInrlRhOnOWlMvQjSc+v
TgHxSMlcK6nATO8/N+YIx3sd6jKrPANZ34VEe/ydlj4AWOtxJKRo5ViIEzy/v2cMPMI0kHllPVp0
VzZpErXvtJdG2k91MhTMoF5TmcafPZolo/5H3oiGRq06h1t87qFqAl0aIvYqI0d27jVBqLGjsjZO
n+JjAWwVBYjDn1TCmit9I58ClvW980Qo7/PqgD1p5h1PZN2dOXOWqYMxMOz1mxbbMBcxKg8gT789
k1rHnbhAKjYjYJlOegoauyXRLyulfHAVsTtMn6b0Z1rcMnWZAnLs8E8cNB+MUrjvCPxYNDnf6/SD
Z9lJYJhn/656GZ+M86y+rzioi/yuBA+2EKVQmypcUGko9em21HLMFfd4Q4vUEbEP/VNDjRninvUs
15TirL/ckx1jzyeDNYBuEJi23UgBD8Jf68DYw9ofzqHK16B1IW/5YlbTuQ+Y6Jq8KFUuFQcOiI2a
JvbTwc8N8Eo/ae/5s95xF0ky+CmugH3yGFpl5sWlHMJasJArynfJYXKS761Fa1F0TsX+5arPWuRo
Hsz0nxOmwidk/a7MtVmn9zNoRiVMg71ftYVlALfgFG/KyApyusmrKlyfpwmdXj1kA96ToKvuRA8a
pmdbmwerltHPU3pwiJTWhBCw0FofkzZNtnKkj8PKJ478EQ8J19IYwTNB9Du3ZdfFuIu5Fpezrq6F
0+G2GyT5IkM02UMFJ6AqpvZPuaQHp66J2Tw9lzTInaQPGEqB7jvhTAoU8VH9loKekvefP8nxLtGU
F5Saj4cB3Kz1N/n3jigbU6SECgp6oaw2jiZEWtX2BMnffVQH42VE/4NdQpBRFS9HwiKIMMYRn3fw
IXwae/veSZqpMWuM3NI0sLIz6gBTDdkE5ll5xGbMtI5fM2NtrxHO4wXQWHJqYNDdmSOqs1k0SWqU
LZkWe/Dikyf9/prjIyLmb1y4cgPIrTMr5lLi9PevChn/oiAjApSdeljCo7zb/GPcwSTF3fNcnIK0
jsAKKuydizadagwAKRGigNYkibYc5dxobZdna9xeO6rgyYk/3nf6XaVr56XNz8QAR/rW1H8qaetU
PoQjv6M9n/AmqEivtK0a9JRbQpkamAxQyneEF/kqoZyxClsWEq6Yx4xW1uaVDOD+h9D0BJ8sJFux
yz7OBSEQLAuFrt7EpMZYA9KvF3JBujuzF/QiLeu83TJocowXpASZSqDnzkgJ+DbfitwjMMmV/krK
/3Aa66xDyhmGilZHuggBDEerNtQC+GV6XcHpc0K55b4TV13YViHOFmgZEWnWaalwFz/vQ7p49cUp
vZyX5BSETd8gGzYqrff5EEdK3UIk96i561M0DR5cMC5RonOiE43ng7AqXKOboq77WzgsoJzq3Nn/
sRFXLQ0jSlgm5E2NKAnQFBuebijv9i6nH4ESYKtDlbaaScduyM4aIEnge8UycEaeW/ard4HJN5Ne
KjFvPXCGEtiFnnNfOmslZglNojXzrmaBu+JHtAVWXoNYeRVoCvMaSFv7393QKT0NVwo2emElKq7u
blLCWyUL0LX5UiszWrbJ5ociF2aeyTDlmg2ytGfW/NBMjKGBOEXQrHDQgEXmkvXgEjAia496K+Ik
/xo3S811vV+gB7110GYifuaEwVPRe9dTBDMXWzDmJryW6e2KuU3PZhozGue02xfXawpwzvwFZf56
ubRR4LlewOSNUiDTYYS/d7sE4ZvtCnzJMy3vJj26i14KENeVY+HkbScvKuKLtn92+mxEtSVr9qSA
aYFABlXxuQcNTxtMrAtazU+nIFfIDWcHW2Bgvm1tFEIzozkVZcNLyWITgsDyfejGJOfFtcPwcYRW
XevfyuJiSLwPdWbI6550Vs91op7D/vBMi1bcc2vvybYmL4woHuxlv8k/SyDcjE0iik5J2ZWqELKX
T789mmqhUQUUSMLvt5/kX/AZGQVxZDR/L7IX8uxSjZE0X+Sg2p9rENstbxnm9exIKx67FmBi2pyR
ROcdlETdDPzkPsihUVd8oUP7LCQMVEjcVurfLFSO1NV04Ljt+AThd+ZGF7KK4AlTFga6hVTyu9L5
O28MuHZMPmyeBoypurM1ElKla3McIcvp0ZD/u2MUtHAr9kgyNI2qzwKKrnbmcGcJrzKZK3pnnRt9
pYx3PnqL2fLu1juf8fmJuRb6J8PIAnZexx40w6vOxCNJZ6ZlE3QSEQ95rtdVhB8oOe204mG1YB5/
KjOZ2eLfaxEd9XjBF9UV2kcjlooLUB/LHJjpkVggRksxRpQ8CLFxMpyhGVCYui21aArEjLV/A7+T
xWPtobrnQ5kEnyz5qRzFkJhz1B7khXvd+KgA1k4SuBSe3fpBaxQLnwTaKG6tPOOoe7a0Z6rC9JIE
dB0EaFji2glab+k5xHYR8/SR9X4KTntrwwbtirgHDR2XkHEFibxqggVztqWRtrZB38iVwVW2hU2A
vKjV7AIJPvv3afmdm/VnqX8Pt6g+pRJWVhxlqMvPLyL+U0EaetYUgLstez4SVG7ZDCTWWFR+JhyO
IrzTNpVhwXXlyrfcKudPXnhagHtDkyXBbqOV6jDi5U13WMz1qnhW1cBsJZUZgUGQxtT/8Uzta5vo
XNSJJExK/yJJ5qvxpKTHoQVqc4X+Ge3sHFxG6kZOki9202nnFJ3U41wePUiqqijim+gUhs4vjFDw
U//JL5Rz0pGFaUJvZLU9muntVd9tCp0M53NFzMszVeNHkPkwJrQp+9FmD69CZRyEu4vfdzjtKHbP
AChEkh49aUsCkrP6X3ue0mRS1kqkbjSzI7lw9tVBHc0aL6bUxkIdTRJckdTHzzIvUwjj64k2S+oj
kjNYI56rL8qgcLTW7e7AdGuLpg5WWlRKn7YvrVTqm7FEhO7xjQ+wAU4XRDAfkB34YTXQx8Gn00e6
gUHYHCZmD7y8vZDanZf7Oz+RZDj7KoAmyiVhHX2PE4CM7/TFtB4Jn+J6qB9YlNLsTlU8ZBsdT/8B
zqDT7AZIdTdTR08y7WIKbsPNqJ4yJwAw+gXGPz8Z2nuF9C4ALw14Y0bq+ifrM9v+89o+VjuzGNlx
3Q5yC/E+lZVuE7WkEZCgrhym8BJGA0LFr2aaD+qBVFnaK7gLmYlC0Z9wwczLbzwND3FmoB69gmhL
t4s7qMy2HEnTL4fVix6sPfmEuGEKbv5XDloCJ88LAeNIbQsaggGpdhkY3RR9qWPH/0rk60UMr4zl
oN2rb/ydikHYy1ini3I+NY9lNSpPbPLW9JS7PU9DAqW2JALjrAQ9SvSrUUW9DkG5kaxpo3Fj8Kfb
ddAo76tu9XhbL7Fl9SS/6ad9R2HCJKYnOAh/AfqSOsmOLBcevlTpKnemQGVbz4hCvVdCX58mrCam
TFdM7390GhaOjPBs3MQ5N6TgY6u+uEAkhGs1FSuUMtzahux3aZopeZOE9ORge5k75TT16BvJIf5B
CqZFR6cTviTWXaFUVRyZjVkL83Hbl2CxxvoMiJJvDSHZN+XdNDNJfLyHTtSKVOPcxNTZRuJF7KQo
PvVxReGANSBiy0qy3vWdLgLlKWFM8DDrdBzE1+HVIyKSMSD3pbP/8dcdKRC8xWj9vcA0Yv0qaYhn
YUbZvh0Tl16J20ovWZwAlD1ePt0AW12Upi0r7c8/z4z1xVaOWyXryxluX1jykZmG+o5jx1ZSYh2t
sTawWo6gQOe6IWeWi3owsyyLlxSDHcUborLuuJslI1OF+UqCJkb1SmZpiBWRR1Qs3pJZjKJ0Uyb5
+iEQKshmCunGLd34PnXWJ2uFPvuQsl3Verv7d0knshTyvYMS35wwlaYRuaR5MngN9JbiwRVF7knH
4HoQ+JbhqVMNPFemUW6x2yKPKQDcsODMdXNTZfE7FMPEoQaMp0UmqIGZFKEt8MU+85OeZ03eYINr
+ahJy/D90IvkHQDFtVzlz/ew1Irc25YHm4IfIsAmQ3NZEIMYn8NrHGI2eTIGSshnq328QB9vLJhI
6hLgepEpgc/Mz5limdm+1d6wqw4nG41Y8T6La+BwatXsVcWIxl4tRY8OriCil4a30AbjQ3rc+jYw
boAdfmAicH5JscUw/HxYQArp81pr8Edy2YmKxbm7aaSoUp1Rpcm0U4keWinBwlXJvsM6bwCPFovz
P8E/EeM9a1dRE7ujM5CtX0s7ZqxZ9mzU/go8QYmfIvPgphj41vu4nA7Om/IkAtWzZW5kzPoJ5WML
+jrSsCYNznxYBYbxPkw3Fy+MZkLze+IsktCKSwDyf3XNs8qTMINOHnoZK1tZYlG4eVswsKXkdCpy
vjZfsYwVjYPO1lTWaqALtuu4SstBs3fcNoaGWSgBXDGye6Ah7t7taRG4QM05ClylvXYyVtJ4xf1+
XWfTrt9gWXXpdS8j8LLcOKfB7bP378s/7dGzpB4C3gOjm3EkECX41/cQFWU/F8Cvskuha5r2xUSe
MP+h69i6yhvemUY9ajbg7Ab9w+NMguCXXwiATBOpRQweKDKzMag1raOI8bXLEWP6/Mk7qclaMl0K
NWpn3zdH8/3XxyW9UD80mTHUOQtFrwElYFjw6VgqXzEh1zeZ1r1H77B+bJ3El8S3eciOXr8TnOex
A2qDM939+zofoeiAI17x6E5iXH8tTa6ThZz3VdAF+YMbUAJWrP9u+a1WnjqBMD2RHIn8Avut9Qt3
fZ6gAyIXLYZ8qbQk5oXSFp9I8oJFo+HTPWwOft6Iyq9Q9+rjYgxn9sa5quB3ykGj3qwbKlyUOfTL
H2oNJq8iAgj1cUIO6cwUwfS+enSltvpjNLp7ZKHVZVSwRi/+eWdzINJRL6Q14sOdsnf+ihXRs6zo
edH8efsCuH1dXqCjohDE2Aag0ebPoRyrm4UaLqbXmdiHvvUXEFVQYAGjWzOCwPNrhf/rBPYrlpQ0
rfhzOnysl1NiN2Tx7G12u3e97NWKFzuTyNt8AVpS+0CrvSMz9LnzmWktTnfSodEKO1F/2R1UA3v1
BVqaNDFMIwSjRzVSLKbPWh025Re6NCCsesTxebHURX2Ba1eQMM9eMkq90HmlQFA3mSePC1MF/HwW
IIpi0uSmaYcpfZPZNKVooHsvLomHx2/1Y3cy791hwfldAcgwn9D9vln64tjnBHfbaSIIN8ht/nkE
MlqA9sGKLDJPN8i/KlcnDxqzboGKgL8QRzc9wncJbSnyGlBAraK+zXbTfD5s4b4HjxcnbWt9IN7o
iZ61mLPzlUx4/4y7bD5UvA4VZtN1ZWQjHjvWsVytxdTsmpQZrLynRiAHHWvLkDIEZEqQi/IYFjW8
yS2ZJ+b8S/HiGRvXQIes8MER1vz8cckVjnhvzyhst9+PtYNAdlWhBBRjWTqMjp0WQd4NK5THa7Yp
M8ja//uacIzwh1T/hE1HG8M2JxTqa6q9x7Z6I1BCoAMj0RNERWlqfvPkBbB1EQfvHKZPScO8jrTe
yi+cKDWktXM0DO+yUpwHs3WM8SlKpO0cZ8pp/SzQAQR6+Z6OwR1uAlVPLmcKOb2BonYONQx5iOcL
4fhm0lrYxYfFsHVfwRHmVcCRTa3t10JcWFLxbHuWgLdwP+GTskKyum2S/PIU4e8JXqMBbc3msOSQ
xlStlVjuZwmVeyX6QL7Bzsi4qlySgh/ChuaUowQJdOASXGCf2Ye8s8NPeah8aBofSPx9gpxT+FQm
ANlpGdghbE+OUCxz/aUMjtkQhdRMyCB2QdPIoHjFuri7y35O3RV2zup1yKQ6eZ2gzfNYAEoJFmLa
Qzsv0h498MR+2+u3D0DrmZZTMm1TMZr/FRGtUVTDrImy1ZFFKv2XdaiBO1rrLCYRdSXLWOXOLNld
OOLuYAhsYtkfypIsPkdb7Jv7ZEipg6PstnbJVxw5s5bCNS90bgmvhOhO8tdGFZcAvg2u9OPbZWKz
5KygADJsEj7TcbojKu8BAaArS8f9Brv/ZcimnZ7UxTt98gPm4hum3DSEe/IVMOpOVXOggc86Hmsi
ghQUQe/HE9omQ1S+M8FV06+VBVj91cBxIQfGAaR7Y0lSgNu0DvhQnMHGlMqnAcoR3mp3YLdCej2M
cjsX54s6IhqU3MoiJR3ozlxkndnJWFdYJtv7KphpFjG/3agYXGbtH0uW5ruYq1O+IPgavya2wBO+
7DcHPuafO452BE8Phk787RQ96bQEt93FGELA5MOs3gnkc0Onf9MWw5TnSnot2Zzq0mlqhVg0HSsB
gUd0N8AcmwmSVXmSGDRYuXQZZ1GGAOAJvLLORP1/bBtZPC44iF51W471vV3V4NYMc59ab0PfsdVx
rOKIFA/hYbsrCJRUHTUhmPjO4OjNiy2C6osJkuWb0S7cLCz++DMwCwhkxrkh3pCMnudongcx5pk5
MdXyU/JfTHTj3L8B8T7/KVL+zJ5tiEIqVfX0RRDUHBCzMCul+NPEG1RfspJ1J1TeuleWMkQXKSxj
JIb9IXw1CTkSXEIWz+i8UPUS5LgnMA8DL+Ws3f3cr2fnRmQTQMiVDIfiQTRmmdZjSEExQ4w/N6Lw
1jfjlU3LHAOD6zkCBb97hWCLbK8TX2fLp7FpVqMNYW02smQX0Lxljd8w665nfzsLyQJHqTyMhXsj
07kkAYu6k97mUWetebv4kpJl0qFq2dyizdGDz4ztTOtlBK65c1YJtufCvxcgCXRqDo0FFQKfvyXY
mEoGftgSRjldikNn565cCRUpQembHDUfJsXr7uRfate64bEJXq7/Wrt39zCA6MpXrV9VeGqNcfKq
q/EZOIea7/q9nWZZIyFIHtBWCIYG9M2wY4bZRkiKi6nhHSgBSYwcgk6PgrR3aLlwNHlZaq4Qb1ki
qrOGVgzHQlEgII4L67ZiwmFqKYbY/hMAarGhuba5Wyyegy7d4EnvO9Q1oTZCq7hlRkY/5FFMyBd+
P9PYjM8CEG236+3RaY/pyip6NfpTemfoBmnm4rVavUwIw1zaR4ne23mRrY+ztlALfuLTYkQgtzmN
yCTWv+o5FD83A/ofL3jnnHGHZuUJHMPyf83/MD04kmCu1ZhMBwBp0bpHxT75xm+jSmVjT3oyCGRG
CZCuXkRCAxM4Is5fu8hpUrm1B8Njj9EtH97M1GUABaNAOFzt8jhQHHAbjRx4AK0nbAsVqbdBY0EW
WYjuLfZsrAIo0MEedpfY1vqz6DIdJC+X3So9yq+l358Hf0MnzhRAg0bzLnItpsqv+43SKm/z2qqE
VxmF8KEdhJVKQ0b0b3C/nrRh13BV5KBh5QZD0yMJJseBFa7CFQCmQiPvYlOgUFcS6Tg0QoiOttQP
A64L9ywWhnykguiGMU7ELAB9tCaSB/yheM9WqeqXzkWkFK5lPrwVe/i7Xox2fy5OdyNwXSCSy2VX
zT1jRYZi7nWCHwurqg2G+1gr0KxE3OkXrMtSKBacSK+HNswaWWrkr8yf9uyhLSnBc9yAUTkHgZW6
K+oHev9dqeMLW91jC3ldgQkIBZnRvuX7cx0GaX1vZzCR7I8TzQzAPv/X86GMcUy26soUvwC/9eK2
43scGoEALkWrZ5CYh+tWxJSgonqBY57clItHw1oGsFr/lW9rzdtYytANKoR8+IQStLTSviPBDGE6
FUgTogP1x3L3YhWwIOacza7zu54oPR1hz9ccaNNCQJ5kYG8QL7fa5ND1kokX1cfKzbU9YuOr2bBD
+CDKSNVUm64OPPyKpYF3Ssx/iWq8mstJC3ogiq7M/X3pBSiUh63R5YrSX5O00ay3mZhZOMzadb0k
kmCat4SWikp9ZVf2+ku//L2kyLq/aQ6dCZ/NRTCS7+Q8DcrWRPsCCtcC8I0wYSSe+OT6vSglVutf
ZtcJkF82i5lUr9R8VMyYTHqXQxz7gJSnKNhVQne23ceUHTzjmoW1u9MoGkbbR1oQktfX2mI73f4p
hCjsp9CDsT2pum1W8itZZAxZK41lQ8xHzGTZndOSdvixfhCUHYpKqo7IdSX7lK0VrTuuCy63Cpu9
gDH+mKC6WlEg7QsomlmvAGG6SyP+9pHqTbigIy6xLqJrknBmW7ZawoAjJpv5IvN7Y6vtoY7kvwfu
OzAZ+PZvxdyHGD+5isiha8di3K72Yy6XGX2Byy1A3tiyMhEvj2vkVji32+1w9OVRb2K5JTGXk6SX
lLPrh9xgmC1hdOv30T9Fzelo6a+pioV7vdQkV+d333naKiEv5WO+pimyxXrZGrjjZ/UVBCqIYoVn
hlJKtzewfyL2H+dMBgTS/EWYPgcFtLaCTP7EvusSdgQx2iqghKoZ4VDE29Q4csbuhEkg6+cRseDj
W4N9Kr6YTbYQZv3h+85nbWo6hiOlNAy/onVCNSKUX5TMJnEZzBAZYnIaXISsRfLkjsXBYn9u4Ihr
b3oZmVFq57Y0u2Q+KK2IJpywu4IKbpdbeAomBuln/HrkDc1SskkbQD3PcMTp0ZVzcx4HZLCvQxlZ
+ByY4gx8U64HM4lMGI+GN3r2TVVXeAouqSC5MZt2NvLMgsNIUJteQVM7fxe79RhjmqLKt5wYB0v/
NebssEIIK6g2uku9Mp+WPYmM1gSM1IAT5/Yz9aI2mZt4K6+ShlwgSIa11LCRWRff4lQxdlqbT24f
S/in158VswqIBeGDPQ/T/4eS+Bd6KxRnPk996+79OiePX4nlMdem1isU1i4xWjHfLq2WEkKPv6bc
4CN/4XelDwuHZNfJhp7umwdAc7vuO3I7v0Ci+TmcSgYyTqKLqI86E6qhj2p7IGi6CGU4ifPW1Kyi
1c+sJ2ndAZZ5JKgAeBJBOuyyZdlZn2nHXdyck0TpKSDpZ+ZQT3kHJQUkeFzXj4zKyXg1WXSXC8HY
FTXT2TpkgQpOWA4WhDTasiDl7sUvRLuxj+OqdIwzwxy1IPbovw23P+LmJiKuB9JRocMxKW2ObhQ2
m2rUZFKlgIbjIz9KtMQdv9p2q5UrcUS39Q3c44Be8hgnglPg+dH8wAcCWrmjgFZAj7gEYYjfeQwC
zIRdu5qr3WT15U1jMcUiGJgVwL3zfezUl7N30yNTonJoDIsnzKZBQEeAY5bjZjBxW7VpOWxMPHja
98svgbAgCwwLuFxeQBvjLKYJOdMOMXYczDAz4SKMLJI3aWgln7HAaPb0nSSQVgNAEFA9Lm7OYXNg
55Gap+Ejtd6nWLl8izBuNDNZLQaJMYOUCGNDiHbQLUlBOxMSpLqgbudlHKuNngAPINtgFQAvklCc
LbS6tg+i44n9BoxZDknx6lhpRJIzVQPTyjKi84ZPFmu+RROBl1inFoe8s8fmP1qF1iZs8oIfAIP5
4F8sMuWEpQ8IjswKhFX0gfnLD/jAB0jMqstiaxkQsIf/BIJD92M3VDKGtYTZMT5yNV1rhSkt5C9a
h7iDMh0uIdzik3BPugcpGwR4xL0LT2OUbpZHVoMBmXY7VWP2ZPAYlsg9YP5tJqiwqU31o9mSE3cM
EWbmNbIqV7B0GGuO44aEOzZWYwIu/GxECVwT5LaQeJGICEAIhZqo77lzGm/Icb+3RwpzP0ty3O9+
cfIGMzDZ4Bxd5//kCqpRkGsGgGKYg9tyVNu/OwUKsaqJWwZnyFP1O9s6RY2nRPZeD4ccvUddCLX4
RTbK4JalReLPuEy942+L3GrM1GaqIgvgtKJBWnhBs8yqsLQTROM1aMyh5o4bOgVAKx8yxSC45MZD
epUuwiINDHrcFdNQwZVKyCdRC8AVc7QvghzmiIPbE8iDQw9S3GNu3MvvwLR02UwJF+SBVIk3DXg+
anBiwvy0+4pdjBm6Aq595sRegO2+Fy/LOd4orjRnAJavqeySrlAzOlXLPMefKA0hYGUzGVfAK2bA
IJAqbkjBagFECp6SC/69wBUgXv/4kDMMGrsp4tc02zpz2SwWhu8YVy/dmqb5y6R0UbDLHbyCPFU+
FecpeYIyNtCC+AWod7kSaN6MG/V6Ji6ivfuDmDCBgDOaVQefTb9R7ubaZAiHOitrAspMLYgcUJeT
PoKXtmzmLW+32Z06VW9bbqeMGWGW+URBletlxKplHL7B19/OuZSfmpsIyXoA6t5MWCkrOjpFi49H
N4ATQwQPUpHAh92A/o0rA/DendsPnvemKs31RnLWxLTKB80GVDQ6wnEjpiBSK4f9xb8lQRQfKYZK
Br46PgiQg5QRivfKfeCwjHoEvhpVHvjv4YcS6aC4D67uZvUH4Wu3KoRFKLh/oMj+mGU75jm3eheP
Nr6UuWG9l58IYqh+xj/BQo1OmmetnR+b21URL1BDUkTcyLochsu0KLU1fQ0B1o5eO6izjhMp6/hg
pKPH7RrsVr7e8+7tUPmTpG3GJZbydvQ+MR+/OVX1oEW7nqMAlgc0zom7fZdtU41KNU/pm0S9JqER
eyyobTDvm/HpRQzSTRw6hGtbACYqNkpx0SgBZnxtjZQdHb7rme25Nls4RCmvJDzvYtiqmWAsEgNQ
nAdYOWg1GYpUkGfd163XU0BTepmgfTJ8zMIh5zQUNM1KuB/rfg2Jd++vu8ETzI20+Aw8ZNvVAclD
wqxSvgJWa7prFqfFu+Ewg3rZGJtlp7WX0wFRruyCi+fZsBnzSM9eJkxk9th2CQpTU08g4tUlXxg+
pP9E/tEkO720sF49GMhh6q0tiUvqaB7bifFKkJVuRUb4WbxNS64a6EcogLo5tpUozhHv71Si93UX
VjjzutGD9Q3JVo+qIZd78kcaDSEFCLpw5g+g/jPNA+dRbcxVADFHagqeMzQ4BZhc9WYpisg0jZ0k
FkMIW52QKJ6wt8QlNHzToo8Q9q13Nz/7h0quoclc+51csTgzuIRp+AmjNRbCp962pjvjQvyyxjpV
XM6WwtdsS8VUK57j7dfL7fOD3Bzpq8riC+yl/PoH0QmcHs5xH3w36xTH1p3se32Hlft2MuLoOZ4w
CTNyvbpvaIaeTjvcNbk/B9VtS6vVM9qebuMy7U+lBrrWy968vosV6lr0ncQM1mTc5gJ5GU6Z70C9
oUyF5rAgAe8Q3FclNQqacyGetlOly1nSDNKPfxFKItdQEEhsNo6RAluoPA8CslnY9wxdlQplo7Vo
k7j3kJG1c6q8UCINfsRuj3OX45XAkFGELI8TmbVrn+VK4ONzqehnx95izL/SjBAMJA8DCnq4QwvO
gu96b4Xz61y75wYKYLIIeEY39a9tzCkOjKSFgxFK3YrXrhuGmcuDNnzTl6jpOzoQQoYfULm6B9uO
V991wooI9ngyiTAQ8i8/zCP45TZaAZ4hzxI0x95Q2ceuROGrIoURT6wVkjKQBpAyYxNM89Ok3FHK
7EyZ5va6XWFfQSbmtrWRL5FOdjYjlI+1llyrZRW0+OhdgqCb9cPMTipgDn8fB51iow8pj6mtkI+A
wXNIBQ8IKrg4agcxW8OiNvA3GCiunCv14Qse1R+irRJ+WspWvC4V4zI/jom/+Coz1Ai9UwPKXRZZ
x5b/km2IZNWnvr0ztbSN7GqOyHzHvyptvEjussXrv4QGEAPb0ZzCledyRKRq0azMmAgIxbceb7fo
WjSScH+afxZ8hOX1fg9ukOIQTMkK8b4auhYmbOuP1Btw8/3+KEZMxtLYp2IQI77GsuM079AGLNdA
P8fsiMdI/Mt8WJ/uyVO+khnyPud/DPLezm5JQKjDC6+2mxHRdT9SaXj/B5dRiVUFBUWzBGC4luGy
N1bTIMr7f2iVyQ2MlIAuZ43XCyMipEPQ9nG9rUNrtc2wv3zki71wFE8ESeeAnzBKRW8mG791HqZn
0XUceguddrukwZrizT513HQBQQHAzR5/Eq/l9cW3PAX+ACG0xInYV2HOF19HSe7LzKPZk1RyEXTW
w2aWmbqlc/Z2YvP8AxNSJrhU231T1ofPeJJ7ioV0GDqxGsv/VSHZSX12mHcZOQe/3jXcArvZiqWA
4oomzezjSr26JMaMy9zNotKrvCEfU7CuOT6SrMRaCDNPHQTBWC4Eqmr8KsIhk85kDZj1dbP/RejG
AFqTTC/BDA0XL6C9PrUPOzvHAyFQr6/7Dg4VDJhCgnVk86LZkesl1o6dOftcaZOAcnHYZ47QWHEA
jgPzVNihnasC2GxKJqwbS6ookrPbtlAOWTdw1Z/2ovPU5iXcdQqahHGpRv7I7mJXzVjsxnqTybGt
DQT2QgoZr67QvfLRB4gbpwZu8h8SReB5EchnP7UnJhuh/t/RKVz8ChTc5eObzx8TaHOEKgE+/dlD
wFgEFTKnzp9MlB3tox6lz8oD3aYjiP3TCyJPySCmkZ7nvYVzufjLzNYyWEg64tiBAfIp7nWya5ST
Y2fGDzXu1pehXqmQMhz6HA0tkMTkErN/B+Irs9HKXgn1fp0/abY9Kl2/AIlewOsZbEAcy85YCVgy
Wxs40XwxjvxlEDhnSVDn/h02QeM5ttvMYcPMiRp66CqtxTn9wmEvu2lDFP/poZvNFJzIoUUONGTV
hKMUffJQ6PYRJJ1sFLG2Rroc9ZQgaNhIuTGu7zT1dTO+0wp1oORUtxDEDu7RIxoi0ST3Q1gAXuiO
1LkyoNdO9XQl/DiTg4hR1o6FzY6Lj7EcNtbBxQ5VCg0O0q+z074nor232RT5TPK8DhialFGg/zgE
n8JLAtPgmpyc2a961Nh3UlzOAXguBc6dP0jrRjUI3bRKf0K1jvRD/0e75c0Aa9bSF+mnVy8itF9k
KB/4NgS51aF4OlLYDNv/BGGIezeqrormuh0afziRs85kKt3pDdoGzQmWW+mbHr0pb0T5VTdqRe2C
Q1yKzK9C41J7Yh2HWdhrhlWqEt6NVGDMH4ySaYo6nOzcqR/HlEQWhJknkRXRVJjkNsa1C7kiGsH1
esSltRgeIXsUSFNUocT6ACC7qHkWT+At0pnwRe/CCii4t+gJlx/zQmr+2nZ/EMgGgZPDuaTADsTB
OLpQN53i0u08K/UMqzEe/V7J/s4is0ka9ULLPa5Oqvr3TVz09AqnL1YpTVcrGd2EwLlBkWD4UwUq
g44v1iWCYFyGNR3U2xbT2BEUneZnOkopRR3mnVPvlVgH36Jiro1ZfqPNunWHdqj27Z37ZAKQKHvl
eVWuDDqEaTLt//Zh/Q4FZcfFgiL1dysrbvUP3w9i0VdTetHf1zu+c1p/o2LcbKuVBmqWGFHlLDwI
b3dkOHFXlGN07oFvX5fs9UqjHfrc94gE5ygb5/n3eUx6GtEu58Tw4L0Hcte7TgNDF4ECiEOiSxzT
h3f8IMLsA0jqifHAJO2IKRK2zs9Lqk6v/vPuOCOCnluESK++8t+o60oaEpNNBnBjUMFCy08SEQB0
/hnfLh/aJY3TEQYoxY2BrsAz20hGj1JSF08ajuPBYyeXZDYCVhor9qwpO2EUDuawfGP5amhQ9h2J
l5wJ5B4WhvwmYIlkD0o6mSsslcsriC2t24JZ73lCpyRAtlnCF8FRcbKj2uaPd7wXsUTmuI5nn+BC
05u4Mvj8tbCLDspQHCAL1rnK0RmwAPC+BX3fjdistIT6RMiSRw8lgdXlMJerH8ghrPY/HBFMNmEm
9RYGacrxMdxw9wHcZAAoVRbpLg3IlPjTdhAZWMVYgWIlu7hLgjvjY8jC8sgnmcw4jVLhSMotWwH4
1vM9hbUnWN2VHbk/cLBl+3C3DiqG8OMwvCvyu3JVtl1oDHPU37Rov14FqgLfVqdd8WfRwwRAevXl
QmeI7pPFSRPjniBj08s+kkffzHlfs+QUbSq7EAr6aN9/yrXIMuJwXOq0P1mG2Aae+BPBOWhEfAOE
Qo3e53iyzNE4vrxACJQjjfoBubReejPB9wkv7pVx2INRKtYMxLWw14hZ9XRSq0yKmEqCkuf5RS6G
7EDSV1YQf8Qg7TBHPQ4rpqmhzs6Fx+FWFAuyI3LHf35MLj/VcXDK2njGDHFsnOH8VRcybbFIp2Va
bHDjNMKMM7Ds0YyBo1DwMH34y3YTsfhhafxcFdJ+zUyjWjuhrydWaYNRL2lVH4HOAvzHowAv1LEY
VvvuixgWCDlw/oJuzVWrAHZPiCcDOHQfK5JRLo4KuoMJi4KM13yJrlgqAMmbayMsZJvqV7xl1qsR
ZLnCgoQJrq5Afn4tILS9Uy42ysk6SW01Jy8up3zlmG+q2H8CCiUqxY6rXcKBzQDZUPERY4uGTCY6
Y+LVTM/HoIW58XBSx/m78/ftgSHA15JSkPPabQlXrnanu/GSLfLHSPgrrHJsHx1YouKTRrc48Czr
GMWCuCIKoNOzarFImz0IhKR/tV1GKFUPLXr8wv8Vp1uZf0b0GJ1geq72c9g1guD1DTAZ5ivBhsXf
cSHSksvMyLj+lu0BiLPwxByfVdfhNcepadDDnc2hNz/dWFjlLKK8dhXQQAAOA2I5CJ0dHZkMy3d2
bP1RPN7Is14KxHSX9M4X6l+JZQTfMYWFsZjcGKhNU4o8B2+Ww1HIbbJgYwSShw/jjEi8w2Jj62vA
GQDHMwGhHkhYtouBjemAj5YutL+usgfj4t6g/85voy3CmoT1iN29uA31GwVdu0sod3Ijc0yOjOnt
i8Kct/bPDmlxz/p6fssfTnqjjgQdiZeW5BqGIdekWHde2CTdV3dilCCI/fiaq6aybz9tsDkhbHaL
lMVQVDG0HdiHEAgfpaC8UmP/5MgYYE6bb0vR08nArVB/PV0vYqMV51EONERvjx/m07QdyzOx4K55
jVU3aTY/zwkP8uuwvc7rjq+D7bRAzJvIrwnHdS+z9uQXymJT+IC5dHUfnAAxNXOKvVPAkVn8iodP
LbhPyfzydp+uthIb1pouXpioSIZpCshpFjEgmvQfO3BiIQsPFYjBeUXQlefgwnWH0IQFTzrW5fMl
wDySn/797KoBAkNWhO97t2SPgLSpvh8/vzjtZd0wQu0Z34kxvLplr/8gwpptug4uqtGYhEy892Xl
RvhRBblHAs5XlmIfHPlfivXuHKDdPzoLGf/okR7DAJUcBYgS7cXUxDC7YRw+HiWZ8VF1boqfa4/q
KdGOkHjPQGto9hUoa/+Xau1BvJRs5Xu0amRr6mEDm61w3qgpCHQmDREMevyixqQTIUHZWh0EcTLS
FlBGI98iegfLhJeGqo20zWKJHRPZ4uIt6nxE11wY0ju7qrp2VI/8MBloSuwYJxzmeQeaLX04dac+
qSg96eAzeV03wqWX4whkvXYdZCiEvgmOtUOMW6uyHHps1WfeTBKbeTvyQMI9sAxtLVungixfuDSp
0HlstXbyJM+TH1X+wwnq6cAiCxtHynyDiMzjbeZKn7NKN174ooLB7WA6SjLbG2NJKLsZo/EFPkSB
TOTq8cXa6O2beQ7yzLtkK03hMbDpHiUCYm+0L/zke0Kzc1C3Ks8kC+2NHPvtMTYgamMQRVBfesl8
zHknlGZ/WV2dGaJJEgmh66RX+4fce/CHgBpl1XMDXc6CccH3cLi/QUkesnxkyihbIzWvV5V/WM9N
GkTKquoPEpR9YsKcHlvX8ufYwf8dtJYwmoINvx6pse+eWWr8B/avGbjCsBHD2l8YHXR8otLHUXnn
tTOJI2B1A5s6IW2CdWOLAfPHa4GIrYLk9vTf+bhX7fWdLqVc1RgxR7fYOKdlen+3yrsim29bcAMq
lUJYRYJQclZcjoVIoKOraGda3LSX4IsBVEFZGZwfkoUZIhViS2iWe9y7GoBTdFI+MadxE5BAFP7H
ntE9pRd4D30FqxOsMVRaXTkYaYiCvbUoLn2KP57k5kDjM4eZKxMNzppJ/xVdhSmdnk9IHMBTaxqn
mJ7zYgpY94RkgiP/xfSmj9L97YWW3LGMu7wAOplM+PQgzWvCGu+Xt3IbKawfWL27wX5hXO5vekQa
5qakd3Ib73PPqt9YA3ZuvfGoDSpEotW0y1c/i8kv8r9nr2+waExZtuVVDuBclaTBiDGiCepyCNE6
tNodJrOoEWQ9S7ceYRWD2KsS1SCDcV1jEobVKxuUJA9MyJAw6TDzImJdpK+WnljGv+aK1N9mKUoC
8VbdWW2v05KhAJD8ukYHNpydMgggN3MkgeS3J2sr3IWv/YC6LPjytbVxh5EZ3SQyPDN72+SYa7DB
kLPn77oeaA25ljuSTpgUJ9cKWa+B0K/2o3qRy8W1kqDM96bfRw/6LW8M1UrFzn9yS4k0GTBX8Df8
oNP3AJ3gzNHs35BlpDCKpozWoqSNiL2jzL4TEwrH2l1ZtI1oYxLbh9OroIa6Dlg5OfthL42TlbLD
bAmKZfsGU86JVqoaIU3ACizjw4lH+7Er9eZFGWVIf+DXd+NAKF2EuBi7OnNVF5dthqXP8yNsvb+3
gjno1EXRItxTQtxbujEko544ctsi0GV8RrVvIiNWW6kiZcgDsV30kFlwQKxQSP6agxEQsUB5kUG2
TO/InQVLDPyHDNqYJdpexXB7ncusjbNjFxY3JkDJJ4zGkr3+GUi8kbmt+YoTFQ6ieICoX9RJivby
d9Ek7jagmjYymaer3IVhQIDSCJsOLBQXDEBwWOT/M6t8zcE7HnwXTTqfhQdSi9SqsC+xQPBFsC7Z
iSi6p2lUHldWsZpJaDHgB6ntBKoi7Uqi/fQpBdGX1Jz4/ru871kCKyadpyw8VGZLU/uczEeKKvE/
Xly/0ELVubsDhYZ4eu7ye52mOyck/lJcTmMLRVTyw9Rp7o7sjVP3+tQAysmzzrzyYdwaWrX9dlgY
n1fCJJvawV2i9MLpnResYdPs8ot5n2oiVPTB8mBUUyXDvJ77c9wG5NCbelVimPJTy1ptNtvh9s63
LiH2TJ8fjS9RYroshodSXoK0m/uOjHSZiDY3btpeu3yO7O9U7V8snlwc4A3q1k+168jpzMCB6Umh
e1Q9DQzhi5VX/c/+VxsrQTpW/I3xjdGUZxCotwVUDHGz64YhY6DGCm3JdLrJyCCCR67xbJct51VO
3GFwmJe6GkUYoZfJWj1B+Lf2fpFY2J0NxfPVl7ANRqKIKoVOiZ7IwkyhPzpsgpZrab1iKBj+6rXI
u6JsQKTwCMrQlX7MnMDnPdLUXYO4HjPYyXuChjkeeWYgiQjn03ddOjHQrqzz8yA2782Aau2/8T6F
VrJUjasRRvkeNtuhWVQDFyaqYwGjHy8jS2ppgSi+AcXp29LHXHXGJsl18qrm0FrKUaS7KLNdamEo
XWvJADq90MqJAbnTe6T6rMeB+iNnzDOBS7ZKnJFPOzmxh0SC+XaqXmkgWc5nxZe0ZvMhzGoFwm31
lw5aAUpjFcMQ1itqsgjOsodkr/HOKMnnKLr7vbZEDkPwfArxU8K1DDnDtHrruvAP9D/pHqZIINBH
6W6PvBsjTyPAgE/+UM4B+IRHok6dm+QjGkSthXZBzX6Z0rxuKXHIU6BzxOg7zr/S7W2HRWc3MZrq
mEjlDFpc3qXWtkzk3oytds97CUYmTVNYINMf6gzzu7NDnJSyxERn4cELQNMagwyk8BYA8IVPxtrF
NNR7MAJm/Bkcq3pO/Rja7KZlXlJi9GaO0iXjkJmD7VJcbnG+yV0PLnbsNM1mX1rNyMrdEnWMjHjM
EQLL+ATB3bjRVcdoYuY10UnmJidU/jIRAy8nJiYdxXuuLASZPhO34fmzIAU0LL+b4EIN654jCuAG
gKdVJ5ol3S4M0wAY8RlxkpbH5Roomtg6iECYxgLYiDWlNQ2mowUctPBSRd5FKBjJF7fGxtBxGY4f
pP6Gcpt3M7JaisTH2Q3BCS5qbb7D7N4vBDLPH0df02jMb3NRsNWdp2um7/zg3TohWpNCxSjTa2gN
Cg/Du+uNJHlgHT4P2r0RflQokQMTL/pm+HWtdD8KGz5d0X8lqdnrEQI8LPqY+p4CvNjCnuKWH2LP
OFcSbkPUFxp5PifR0vFGR6YC4cduyX1e00l/Zdpj8qDkREANxUcgGYBHiCt+1WExcewStP3QwXWf
bBd1503EJ7b7BY6tBNqLe6fSiW+66KNZsyOr/SMOx8eUL9gRVvGEff1Wtn58Tg8qAgzyQaC96mD6
CmmxubUZnqCsfeR8RNALp7BlfzaTlgSpPeEur8d27DqTS1Rn0YJQM0IQPGmurVPY3FjEuKJhGqih
RMSKnw+YciNrrpCzFmqe5g1E9FBx/6EOjA5gpLlObf2qr3T/FC/gzDWIjn44zAfyzX2WM/UyCbhq
rWtwhMgsiepsO/LuksBe4TbZo/zH7J5nCr0FR41m9D7JBhQE81WtfHizTdKHiLb6zhzdSbYMGHhc
pQYcgIlhU7ksxye1rRSaKr05UHXzjZA5MwZSxl2JmiNBKHeA4Tf8iOak57KAFp5A2BJz3EVhr6dz
Lp58cuduFI+XjmEfJ9f9DSA3k+EfQU4qMrx9wNFcz7tsEBE7fB6XkpgQcgA/KICB/uA1DbDQmVkO
nlcbVTPa2AMwtM/RLzt+28YHXf5u7Oaufwt+GtHO4XPjbbijD1biFa2PGepGVxEoGw/5XAdkanZJ
dMosD78zTanwi9JrbKt7LWr2SHIYVJcVZoP/LymIexfYXFsSAPQxXxxZHXN3yA3OCYuHTHJs4vjM
auxipVqQMe3/wqtGcp0KVMdaJvHcfBpzarDOuHKFIJWqRSdhw4VDPOZZyjHfjNg6idk7RIV6pUni
RmMeMjpSU1oeDYbvLbI7wzc5bVjXnYpQky90b2KczwtTZxdjIA1B3IJAbo0a2aFEalGpt77NAHxx
Us7xI8MLTbGEB5LO0HdR43k6HZka/51k9ycFjZSJ1b6J0xA1K+zsV/HE2Q7TOfcKyPXn4KplQ4/c
7e2Bb67B/al7BD4U6aUpCkVjYLIlVFs5qoWwD4pKtA3P1LDBqUakAwKq7AneiJJlYEo/MOyz1ODN
ef9ts2t6pim6aUQrZvMRMXV0K75P2hXFsNM/JXyjl0zA8FHMRgtCz3a/CCm5NWuHED+JHkcSUcto
F+yqR3/Hfo0j63HhJndESQvIbWWOHAGt52OPDzYOwU31mmA05/CFJDjyFTAESTqtFCg/d+lA3zp3
kw/SMQfKwqNghAyanEAwEPEdr3GGIjKyQWiC/FY5UdCTIb5jtvFq1hwb23YLFUx6uXKxdyc/YB+x
q3mW7skKFvUlg8p+y6cfphHr0nqwGZ1KLiLoAkSmItrOJ5z//UHV7uo/dr8PQSngPITa4w0HRvzX
HnfT8HzLePB6I4wrc/5JMZPagIJi7vZKjWaMDE67wd/UUbnZx8nI0+6lA89TSNLSc3T+5EUo1Ns0
s/HIBp2QxUnx31pm0lTQKO/tjMCSERmSVTp8m2fEgXL81u6iTtvuCXfpv/6ABg6RiGpF4RrC62FW
v/Y/YJP3L2A64JXk0rSD8i/6xHnzxoqNC+XD3dGPNDTOueTqEhpj8eNJ3D4v2g3EP0V71NlfWXmA
ctCZlb5jv8pVI2GNER/JSANNC888lIq90dlyQZgTept/f5CbMRcmG9X995xhk/P6mXY4THuOlvPb
4Cn7k0VAf3U/ZbFLOINU9jIdWfIni+ORKERgf2GbG5ohuXz1mKPYUDRqhNH1gSN7tOQ4C9CHwQXG
sZM4jaEqNr4oYWj4K2kPT6sR3av3o3lYkvrp0fzuQvFuDyKwpYdwlCT7HO0gcsYsKjuSnfSUoPY4
8IwyI2RuO1WPdLFQXwkgvURlp2ZrTjzghYTgJkj0EUOntyTIXUvPGVfawfdCjoXJgYA9mnP4lQEz
UFvdpsNAkjDTTfnWmlPH4L74dEhFkyCKJHnT+1gJg58dpsrY23vWN0YwUu1PzBw42xo7lwbnJqKy
ierolFDyzLbGWIYSsgDkEquuFJ45x5mkBkWM/ITHwy2AypreM31ZzZtO6lJ6qUkP74mgR2X9a4au
fP4EvDS0MpuDjMvF5zYPgwCFXMA8eQo/9gcdcS/lX63jJ/RRbEH4aui70aj6qbHMrhTwsGNonEVd
0V1Fcb3fAsLsWZVW7dIjDzqoGXDP7VWZbNsmQ0Fb8XC+yF5ZXtgob0Ue8HRK5MOj1DuJxoEWSe/C
ZzuRxNI95bfPgwvK5vS2SYSl8FSXLWAhZQ+YKy3EMG5blsI+4tovIhmhxu8mj0fJwcISGthsDQfe
jI1r1xBhq/2XkarweK9HOE899e6gs0xRhx6b7LBrgoMjJIhCjgVRXlhP6BDwhGPFUr6guHIGAvLZ
nR1AMqhjkrs98n4CpgzW0hYHJKXeKIMcS2IM6glna4MGkXbKTpoQZhiKXfmHHIDBJlnuXDMU4cGS
PEVa3vsrZG5/0Ps1YDL7eceSynR815Sy25QWYzpURkY5+jIcx3ppLp1EbO5vUaqTU3qV0C15I33M
0QPF2Qh/RTzuCs3cWppw0ytna+JRAxeFrdhpWxEW4TV1vGTO3ZW70jI+zy9h7sktyEDQXXLW4wv3
BrIf2hD0He0+XYgoHE92TsmeQx7ZTpjDubSQPJmNvTJm4Uh08Dm7izfqwR3mwiDfrj1otgrrv/eB
HQ82ci6Iu7aNbHKVSj+eHrE+Qm3lzDcrGQPNpNwqsW9LHNTvZNejO6njiRbL/5rXkPBGsEtyX4HL
r8XQLmU900LJcO7hdlW40Pt4pcX7hF+x/b0EQIPCK4b0TbmLH2uq+i8rUyGDF3CmjJLh0wY7+8Se
E7oYF6xhjKGZlPsDZYooC158/IyRWsusly7hQNLY9UB9bY0rvQ12OraGEXfk5T2M1INI44hhpGCF
uwRdF+AjuYHKg+EIGO0I5mtIM5i1z7pP6Eq8Y8SQPQobsfqTnJYW1InB9w8F+HSQNnpQ/p3n4P8z
IjxoiLrEo2non4hUP3EuCRQlNKRa4wStrKfi6Xg5NXJyTm289CX9eWQWAYMFSWwr64efrP7zEC/N
UWqdUSq2Ua3Uzh4pkowM7bxWFd7oCFpeZccunMTMmaQdkbQRb6ZhaiBxLCvrSOLepeZ/anhdBk3n
iBGghqUK1jpaJrE03M7v1Vd6qEz95xfnMyjLTqwt1mjbhZ62G8xPnv4qdSfFWTspLFyvE/RIznkK
cLsIigFBKUNDJyEB+cMT/w+l+ockSKy4U+N5+mj1nt6prpKzE6a/ekOdZ1yWGoWFDBrgpFTCIehW
tmKKMEeN+UEy4N6SKLFYyA9r0mxjMKI1HydyB0/t0h3pmiGkBWqpsPueX63E/09DVZksasJ7lJQa
1BT/6TX39v+3X0LnRnGpD9sCZhCh4JLH1cp32EdFw9eU20m81YpcHaFAIJpvTNHiPo6uEqNeLYZH
oqqcXNqBfDPHfI902AFuN9LJpxVGyx1o4QGfGEGlriHdBuJ7FxyfX1WXzB/RXE2SUl/7SZawA0Vo
HoOxU2fFGJayvYcB45vd+qO2BAdWHmQEoWuQ6Wyi/jsQSPhW+/dTW94Akvurtmugwe9mmmmSWem/
d/Ylbs2TUlN3gJZMp2mnQDidRXHiRRMbsLatN/ZRNXiAtVYajy0EFEp3FZB/Xusl9bOZmCZwEU2o
zHR9ovgIGUHBdngMAKd4kkW25nPb2wOaH1CvAJ94uhVZ6r0+m0dtjzjjYNmZE+WXiZv/dGsf6gL2
XNLXWryVoPEJB7D/WMacj653nPL3iB4RUNtg2k72lnYDRRP+0YoFsZT47oWds8nzHStmp//9Mykp
OWrXyjmyTeQDrSjEtOIvjqfKgYrAwebFT1aNtbKBmdUaXqwV4II8Yqu/nlQNapgcVkIUJjI57dOF
Io0bKGK9Z12wWcc8R4YLVVMcOphvDnjRrJDz1prFC1QCjlqqwCJILtYs1Sh7qDS5EbRVSoILk75K
11juJwt+WsoKeUo5tqa5Sd3JJpGV4dT2+83y32VRjplMteeYCct/yojI+gMdk0dQGRdmKc3UJs7/
NE1A0vkwu6lk9O0RH9nhj5/vJO5TMxdITQGVnsW5bpLS3tKX0JwzlsldGOMdIJw89qicN6ZmtJmf
wTdUUuSQ4KiTZWVmRFO1PX/1T6k+HSg2tTJ2dCFkcrePZ6CFCjykRAHdhS0N0qCuBkGmRYqNgXUs
2xGdbGJg9MXyPeAMkqwBScyRCq69VJ/2NDfsGmOALLhsgQFfGfmfVJzIc61tM1YKCt/GDjWOUFIq
fIZmG8xu7/0RIW6Fs36hIuGbUpaqVneo7E/dTJL2D2uJKyo0FE2wqdCunjtrHMzhO/A7e+tKsnYB
fHyso0Of4FEadrATGXxb8szUphlEWCn11rcMQzvbV10DZnyxtvtCsqGSUdaIntm0GiPmHAXJdvGh
QrxlTFNRzNNRxUpM1ZrsP+WSJuA6nmzvZWIb+3BA6TLMr7IZAN8bec7GrdIgOOU8XldBAVhnOyQI
niM5HIviskxCxL9CoV0smyggv4i0pmPdUtYgvi9qVZELkDZe5+8paSt3hJwKJuKUEG+UgEWfggP9
mYUM8kl/mwHSkD7u/1SlSjOONhBys1gRwX1sNL3nP0mDewtDvPVPTxneUM0Nsuhx3BDxTdVAbnZm
61vI8z04AJYy9Tx3oiEC2ctS6MxFBw8toYS+W/0i/JmpbfM6TfremfIDpAcMHh8J+d2PHVtyyAF/
L0VSIhKGGIAIzpyMKpcHih1i6/1w3hkVHApilFF9zdzld0AHIyMaR7g4XcPWj7nIqf4/Mc/eOG/8
+m1BwGJOwwxptBAyQ3brBDHDx0mfZTTB9Fj4TU4b1Ochwmb6SiRavCLGEp5Dyu4wlD0QtJQM4zcn
37WVdS5hBBKkhB4nwp/4aB3wJ89F8bv1v/kVDV/l2oJgxv02N97Itrzctay3wf2x3bYjVsePePel
fchUNfDMMD9NcQak1bijEcHCc3biguUIesWta8M2Lshm2J/OhJe4Jk+H5l5I/84FS9RXJ7wysalr
6gMLmB8nMS72eC3X02x50co7APze2bAygtToHbeo+BlNKVHMs865dv84r6Q0RZtgxkfWddK2iLoV
/JKnI6FIVTtY5CXWxyU8Ap2l2IhLCKcwx9zEPFP+M3FrJaDXLW6uBeIa+i68E278GOW06952+vPF
Ztn3CtZ3SV5xKs93omBs/+RAQI8OOODekb1ULZipFuIhVq8e5CFoKenxhDb3Hjah99B6ykBGhdEK
I82aGwAOGJt7IIwZsT64i6taFmKaJDdAQvieyc2m0KOahjg19tImUMcILeCgalV+Etb3d5OmWsAr
8BxmMglVHQQxwVDerUamqSbQRNNXFRrSyfsueEoYQ0SeWSV53xokQGWTXkSGhYkntRgAZtV9vM/t
w45H/kKLK3RmS25ZLPwyRcqBi3VKVyS7hafW+1HU7SyB0sAV6fLr+v6/alLHASi/+7flbhBZj1uz
XfMuoMNEd56imSv3rr7rdna50b9lARSHDJ36S+yOzuxL+Aa4lRdhNgTvURUKyxggSVuweY4rlZLS
wTaF92diA5rucubcrNlRz4DD7kAljShKVXijQwxemgIwV0jtZKtQhKwcbhLTBxkqPXwx5E7Ri3ys
EdNNmSYcYG5FSyOX5neQqGTh6gfWq9vRVSpLqqjlEZORfnDmOof7lyowAYLn73PVSoWykYBBqfnU
ZA/mbwrQbkQMcgq6+GJUG0G3hCd05N+6zqzxNWEOFrHbQaHXHP73bBHIHlx/v5WMUWihShnp8BAl
YSzfSl/9ziL/g1v8KuG3Lju9lnw7kcqLKDdegQTevHuaMhdu85V2DYCNVjQmUMCSa0pZh795fqZu
5flFD85mt1IuoLl/MI0mA95LofWCmllOTno2IaXuhJiIhRJ+DPYGQZyWVJUQwiUby4PvfujA/Cd1
RW7H3WeeYsc6QlYyo5Rr4ALkiazhiqQ4N0Da/uG8kRPYCqcL97GtD9PJAT7Q8t0wNaulC7cg9iob
99Pv80uheAs90JoQa11Ywaz9G4zMqckp3J1sw3y51k+k2p5jKG5QTvy4OhTULyS8LJqX02PLX0BJ
0jeRRs9TeWw4mxFXClm2WB3FNxFgBaslmFvhek+e/SRq6dhYE3eZkjqydMduTqikJoXfhn33IChn
mrI8qBko+CgB4ukMOLSsjaDiaX/gRhdzslugRstDhMVxcbC3en9B7b8BxxEGKQLX5oV1E6fH0hch
s0TregBhOoAcRuFuEHs5fXbcmTVYTySuqPCVfauDdkJgXX4zdU/nGjzblSGeFXthgCAz3NZWL1G1
1YangpyXJwrlfb5w5f4nR2S6IUNEP5ZzNqSTl3dZU9sWcGRGbMq+2AEZau5I6V6geRncJIpeMb4i
QnH87Y/Lb/ENmE26fH+5B2fByp4jHOc/KQTEDo3Dvn/tQetSHxKc6VPI7D/ZhgqLWclSWW+xcATa
k1TF/bYPEjzazrSWIMTgRzpv9BsrHtsnkjjI/afeLOnhb/qb64lbPUAMDpawQ9WSGSos4CTBUMZl
o4EbE1LvRhOJsW4ov6MTFw9pAAo/l8I5qz3YlovP8l5WnLJbjYinh/foJrwOciaSKxfzaEhI5ocX
CiqeDi9KKT/o3OeYExBR0K+OeTdXtQY9RNqGzHhtZR15TWSpFzjdmlLob0VwM3GVuNGtgKMmeCgf
68f4R86XMSkzJCFplbV+3jBt32c4mwh2QY67+D1ROJu2+y3o3WeuU0cui8pYBrEHPw2Zc9qu5FVx
Ud1f+wxy1t0KkD1OHOzUFFI4HBR43VVy8HVThsSzZW3dpokJia9s6ttx45Pjei5OlUHDNT1EJP4J
8nZrymxr2LhbTeaCI2cqNRujprqa3ASHrCZUdU8OczhQU3mm2Xf9Pyl78kIvNSdEUx44HzUvRATU
8OH+eRjrIEuVFp65kl9k24oL8TxeQWywYrqWQ4fmjFLBjls0yREQqFibKSUKFmUWFCfv6GdtMWsG
3TIkCApxO2EkTRRZtYVSOKuoGmwV9m0r7/u5x3rgp9R9TmoT2mnUZUhKDIZTkHuKRDQ8X20paqrj
PrO0UGpfGUo5SXV99q6j9qgnhjw2O+3uHtL/Vv+Ipo00qUQRdUV9wJim3sxP8XtR80Y4HAdcZlmh
GvKZMQhj2Zy7Kf38AA9AX6qatUn8TxSo6G4Hcu/+ed8SSrbyD++/HeCrj9yWm/QNh4Gs+1+NdiHs
h9wkg45gk56vnBq00iZrYmXZTKulN1nvCWWMtuhoyB3lvF90yIkLcgsxlkc4Jfmr+lTCGHHNyfJM
DDO4WAwyzm9m6MBKdaka9nDAwcQ48aUzz+NmS3RQjzTQtIWS7PDcSlY7B1UtT7huGQujeXtrJcdt
ehECxNJiuB27CEhQ05m+ETcVBeMux6L2+Uzkn4vXxL5qmKTsVGDEV2T/3E024QrgcXRAcbnqih6B
dMzWXYpb1pnwWbU7+2YSUxhlWbMxt5r99S/8tmAVMcVotjfmz6C3PdzRxCdervGxGedUsMwogBrK
OfhbBUH7BldJ33ll1N/xZ92OdA9I/nD0YFXPPSWa0FNAIYXjHEmEIxeke1kjVxXM6OA41jPFS7SM
VCgyyhAqnaP99UfbaF0jSBl26Pzdl/R910H/kf2z+bQKXD3Xr/pkZ2Gd6AjXh9b3elBeIb9vENhM
s0bN9uE90lQZfbhjI0fnQPLf51338GGCXoBNMI/IOw8m4cNiP+MyxQUnCNTsT2hCe5xTCOoi2Z92
lOBz7Kery976+rKlOjT/T52nYdBiw9L5ZV+OW1J7M4fUojzuxAu5VKuYJsLtE9g4vb/4lQnvySIi
zWCuUYAJgeQrw5ym/X3KCq3LUtWS9NU6TBKDXWyDQhGueJTfyizjzy58us0AJXYzFbcHsAl9wk4d
xUqJL2EbV6ghWZVrzhEldubiP+xdYdyADmENuRghbpsDn7DGfBquV7Vew1DJDGJhBuurPwwtD+cm
9W4oFbqhQfe36VJ4mcytAreeXFhMYckTLzJyxKHM8HwHaxSCMfnH97jxDC9nxEOFnoKLALJrJB8N
lT5JVvfZ/oMwMBlHqxFj103dYEyb7crSizUI7+t7BTUYj9dbObozx+hSyCXAuQ9tWkHYdwGN4Qp1
9EbNVsimILrrb2FSM+25x6Yfl98dhPQc1IklrAhWUiLyGlHNv8XBBuS6yWn22iBQpGwPo0N3PGcq
c7L1uwcwnR3Du8lD+vKOrHHNIrB2Tr0a4q+oCtJmzIoawWA/+hcioydjbZjGYQobZdbjI7taxXG4
t53LZh5ySLSkqCLW37n7c/1LleyDqB5sxa56hAoLmgVr2nORWGghmEB2hlZVmxJhGzDV9GfLqBXZ
1vvgNRKlaS5C8Txf9wnoa9NDu/Ee0RqZVcTJN+LMxtrimZfh4nFs2Krk1G3Nj70zkC3OBF/PEXuL
/kNpuBnxqD+Ba5LjrD37QpNhahgDDQXm6Bi66a1mazJk/s1k325iJGCIeWwGv0euQfkt9dOCtMdl
SAEsbWVOXpV2w5o9a/U2Tq1PML2r1SYXQDMmcuO+SMGYx6UlQ+BhRtywm0MaYPknsIXoC+WOGu5Q
i+XH7XcNtBLOhfySeSpIaFcQJhIgFcKBcIFsbOJcvKIFFqqmnGsDlrHHTmKkElrc22u3Vz3zG8wg
guSri0Eim/j1IectsMV4gf3JBxdE/dGAL5EahOi3KHcLQgY2JDxf073ZzD2cDCoNnF8s5gOL66N7
mX4QFuitZzAkr2DqDWzQN9C2g5l5p/gnS2IuJ1iwgAYHb1IO1dAsf2H0U7DhhnWtpLAdzUUKH/1j
Y73KwzHk0uFMVTgvmT3KyhIsIW3+vkyjanYpOOpMn7T3CTg1IvawXapf6vQTmS8a98izeaMSc26B
iaqm22ydGvKCZKFVpxPBC6LMQo+To/YQchYzten2KO2O6j1cSlunizO7zZB542m1eGUvFFzQ1hOM
0xbq1vrANSWMUOIPTuO/SeysNzGpOqm2ijkvQbL0lrKqFrzJkqq/NqkO5lbEOWkqIdsONmwvm0v7
Mh+Bf7VQNL0oxTe3Cm5kX2Nk38uSuJxigyDJd2sf3hyT9rhu8fj15FIaZ6mo80hgjKNpjA5cY9gA
5W+Er05NnZ7UPK0XIaFyIB1wKSzs8O2q5z3GQ4SDduVs/ZwlfpZ8XFVjvJnJqRrGzkyISygnKoqs
vb7hvt5TisoVkHuNc2qVu/r1887EFn+PKI1k7SlQbcWrrhns1J5dagt//k4650gxM648f6SyF9TQ
RTUJ3x3kG51NTkUvrmvxxqHWN1nkY6QeAF2IiF+Fp7s3OdNpJZMrv+Yik8lr96y3gw2P2N94XVHH
qhHFJ4wgBSxOCGixs19tJJI3v2awmbmzOKxC8VVbb2dK7xL8QHjCQVbcYmTJ/VPr6ahb2jO3FvEU
FsFO/zDxzlafnsRxjsEeN+59lR16KY9i+f3jsK53KuF/2ISKhKAJsi6o4xQmez0G9YfYUTS2SnuX
73IENPq1JtFRjI6Inuk13YGTTAUz11jhpF+1hjhi7mp0H6kMM7IzUi8wjboQGUOxaJV0Qb4/Yi7m
g5x69GE+atxPBtCfoKSa5XQXwunoTJpVWXXo2EofhQPJR/w0criapxgf02WK3O3NC7XqvT2/Huea
bYUQiuDnl2s1MBbaKFt2BiBn59CfvsA6cZsEmrZ0jVGPWelYCkUGA+yFEunRI686JcUc/tC3cvOn
4vq6wcGHtli3UjxW1vJtRuSsthmjxNvBb14pdjqKLkp9HGWNvrytygMvLPfrBQIiYGgbIZOnr88V
XrAvfjaUGQ7oKSiOn7+LSwOYN4flThRBddf5ymIBKa2J05/dWpsnnFHlfhb1BMiofWBFroSyFQg+
5eCIKoq5yT0SheI0E3rU2eEMENdk1PbyTTU8z2ziNGhKEXgyTkJLpqPLI6EwUs+6eKfiUfEqDt6g
qbRbaL1oq2dD9pxG0iKDE2/3PF8qCHnSnRqKJyjrdgzmOclrgXDo31hRJWMvSXg2AUAsN8PLIMCE
fdq+MTybGEuR4s4RPzmwHuJ/TjViB+n9vk5jhz1rmTvS5XDlkP1GN5st/PC5cUsjBTUI4EsNJg7G
1Wif0iFDcY/xlbrOfX3vBOEn+S55K2ZASe94WrrqBZd2o36+Qea4ttFEe6pPb/K3M61JZhhYEcSH
XYMEO0kly4TkFf9IgQ4X9+pq/ywPwISAFI0CKW00+bJ9DQgLUxsolY3gtpLM6cC8CTwWVz+3h4UP
a72VOj5VY31cMm2md3WrmPagQ2czN2tWYuqQhiq/fJfsHxIeHOYa2kH7lKDB8jWwcd2Ec3hjWYET
QzbK44WsIvvlM85PogK3BPr+z+ODOlbTSiFQSVyW7fWNBqe4owGli+rV2X2UM0z8uM69VHIWosCk
A6kU8ovPo+VuRHJBdLoeBjvXN0Jr68XQRQUihfuqYTRdNYPElyBP37jMtOQ4ChydiCCbq+qpsK9A
yPFLMzzKVcSLTrJzKq6PzWIZ0TZyb0FdRnJZOx4Ja2KhZOddAYCqDl4gqnni3rheMoRtYC66y9wp
LlgBV7wubVg2YT2byUj45DsSIkiBFXmivrrgl/bfvwatj1VmG6GSpgzrtttvo1xjE8PD9/L5XFl1
CCgDQtBkQOY4JGoQqNzcEpn5PuhL69xVpmEftyU72pbDCq5D0299HyYITzD+lfxtyYdPmgjffd78
xPPmOcxzK96edNZJwZ1Yz0sAfI0qWdZfZYuw8PlbmHfeSH2txA6Pum0STOx6FKeVsNPzk6fsFcqM
VkuYUe/Vy/NXG19CGgWVzV9LHbVnJZY9gfSjJqNJklgV1hMa2x/vZ+/4SdDNsPm37dPI6QbEBtm2
v07mKh/thqkKbpK7iVkxNSySjUvoatROwNCpC/ZangXbqmEXF/XTWJr8D0Ubew5keeHM8ZdMlEx6
XkvrNU/nJyczgOkkrsMbydMwnRgB1H0Bv8/EmczM3bprVQhfvMfgkKKUyNRgh6aiF6LysqR2h6tp
49w9noslfi9zDBOc5SzUD79r8F5pC65deJVQkOSetfW1tGgcGeyh94aCdoynURJVAoPTSHRta5b/
M2nwq6KOtuHYx++Dez4Rp2+NsPWhTvQWX8dqR5cq051wUR6rdN2gtcOvbE8v8Jaw/7AOD1AETXPk
qapHyTEllRbVU9fWNnaK/LNPE+wZZmNbGh2QNkrwUjt+Mq3tEkLAWQYfq4QuOhSu3+zdevUjadtN
PvBkEJDb3RPqniPio9aexObofrKq9NUZmijigUA6bzyDVztmxytgTabZZLbTR4tVq0on2X2Lh7Pc
Ijqfn+j0mdrMhOwo33sCFvKX3dYkwqsGu9SPzeYgJycRG535kFCyUXs1QXZjJCrly2kMGJqkFnPh
F9epOPud02YwwUkS5XdubEUnqoAiB6ljCnnHyWg5Om5rje1LDkOMxRzm4HOD6wsnXcDXOHE3BPDk
UYByAf9uPn3ZkBb5+QlPK4psG+pmZAPO6Bs0sOZplEjUJxUqfAIkvrFWW4Cftd7vD4IcLDdaRlNN
meCkmlY7OzNS4kB0B4uQgTdY4EySJnROJUuWyxtfZRujWlyn1jb15NHMznBGu0y/JYiyw1yu3/T0
bXxE+/Cn9m/P29EZGmRMCrWwWist/AAFLhQ7vJ/SC86UkYZ+WiIIEw0sAciKAV6TmLj5GvomYixM
U9mxm4hmT8vKN5YGIGMTpxt+vcnA4Rr0sw7pF0lDq2FXsfFoTRS3pQU0H1Lsq1xmU+2p2e5pxpaP
BvGrjU1OOv3sNZ7H8AYiXeFPvhFUoUN/MX0L0Buzj6O/4IS0cNZ1hv9kxKUa7aASrrYdXCJcFFR9
PluaGqFcxnJ6KBwalYwDR1TB1PCQcD2fbC+1cb5Kj0QdqWqAX3vsPLtfY1c5xYjMJwN8zQeOZZvl
Zr4hOczCTwuHtiwWNKe8JBKuf78L//drGX3KGdRqB8GQZtXMSrVlNrSpqpp8au6tNDb9E3+jZR3I
hAL4XXnGNlka9dbN5+C5V3RQbSAQNG4L2YDd2RpupprsywzVANA7xMgvf0Bvw8CSUKSvy3wSWOKQ
zoFSaLhpa8dcIx7jfifFrOjK+V7raKF4E6zkk1RbvVYN1Q6W2kJqVURfn76icr6qWH/e2CHThDu+
KbGpqbH+NU7uYe0ljuew8OAb25Dx/wtbGSexU39ATdA4NcRh4wnwN6npy6dwjIkXhVK64EP6zrUR
FLpr8d7Eg4IBQwhb3sBXAjebvGZh2GMRpt44/vQSqWv/bv/OdYv4ZyzWlkkdkyAzYXaP7ywuK8cT
DM0q0/sjDIJu+mpzxOlwbuhf92rzn56iVlWnhgEgUoA3cuTvxuulkGdX8p1WckNzNT/0R00GRtV/
ivNklIqIqIYPhg+waTLGiFT/8GY1h23omi1MRc8CHheIljdZjoPefs/vnsj0IKmbcoOcuSycyK0j
5lmKZ9gAjC7SUIcf3bbHYV2nGbVXP2nUFTvib8ui4+7u8LFASeI728P6XPFmrD779tcVV57IaWXf
U159LooLa5cHmkNKQBykXWUYP4llM3zLZ1zPNvxdUz91aR0gSU1Qh01SGpEyioEmT1ZyTfr+NmId
XRNp/X6nz/G/ymuzepp5InPhFVTXkIAU4x+J5+RFslplS5X4ixjmLuQ0i7W9mwUUZOrvbQ8FwDbT
OY5QsmoMcuefEgdMgDbcIzL+tohc7bILHkMhtm5ZIgXgvZDx6mkfkyx249ZzZSnAjks7bgDimoMv
z7zJFFe84+3y0aMSN+h/oJbBXb4Iy6/zdTkkIPXLdCGLasYv2W+sOKV2JjnPMaHdVEF/6w2cRXPu
fJ15j3QDlwx4ItClof/+p/PLGOYV2POO2WN7QxkzRhC7TC5dTeTKhUXNc7lxw29ohXrIpVzHY10m
xcpSQGHTdZNkAlwk09ZDt6zCunGlcPQvzH1WL5aGBZpFZroniQtmdGCbMxK78AsJmCTiBy7FVClm
beQNci/PQ6XAd9wKn0MjYlb51otf5PLg9KD1gvSEjTT+oEsERHamvrwvm1QKPG9kfGx+nvMCYJnK
7RHxHLsHsGfhpDW+UzG2PXXaGnVI4n6MV4H+0zToWyLs9QKlmCgGMzwYNzoT+e0QgRdl/xepp9en
phuiGDlle3wWwAY+RkNUxCnTIddnhJxjG25rtaT314sRP+FTkv2peS/6J+6OmjWEaVsA2AgqN8oP
UTyDnPWcNOsvCQEKT2/k3E5JQG40++ecWZjUF9y27d8Y/wc4mhQ7sjZahCNCIZz0dEpcW6F2otSd
4Uu989YmHrsRRz83xawEqmIjqehwtVlPG1Gk77e77WnFOPWzOQ9AHgPPGjDtqZI3Qf9Zzzli+VCD
sB7OOE0qaU5vvaImlCdylW67gugCXN37YBFSPLpwgKGXgZfDzChQKxJdyGL95HSblcgU3uY5SGsY
Bw118fEnMcsCngjIr/di1SC7Kwq7ClDB3e1WcDftdjcEbx8x0iSBCeZzp3rdNfU201KNQLV+ZJkB
xEAhGtgV1Zw4Mf9PufK5jff2vXoU4KO0oYYX0G7KQeLxPzXT5fzbCq8FlCIhd72nd/tO6X4iEhD6
rt0VRPjkOd4bkwZtxeH3YY2OowvtUARSbSns74ZO5oCt6yaY2b32kg+PEpr1wEOARmq84G+EFY/U
ErUZj55KcQjaKS2fPyzET+y/810s67RDkDOUKTHT5lP0ZoRwgULW6vIwwsrTk2r3Mn2YSR3gOaA8
b1QlPv3YV9dJvYcicUCGbrZze3DE+KPAIMNuz8F0/oQp4SgpqQXqTnl3zRACrmRYAlsNTMHW7Bob
GM5X3mWGoWWUfP8UViEKtnFe/TEAc9ucegrk1EdGOJtE2A7oSIY5605D7XM/1G78M9I0bk+lQNce
vwjPiyPIXHOLJaJaI5g/dRPVVe6zlmvOT2WR3du6dWZlZoeO86C/iNbhjNfuXBtYrxDMWeC7T6vh
cQUx4LmwykIo12nZgBbj9/P7hJF9Id0skWlFl4jEu5B/NmLFF5xEzAjIz8sMs4DaOCK+4H9Geot5
Gd+iTN6ZqDumjef6fFVw/cB1nfQ8uMONAqNg8ZR79Yoktoxm496nhcEqta8GwnszPA/7GeDRfjXD
7bEAMt+vKEZ9V1kcJ+vUxKWc89xOK4GcABnAp/4pZLZx3/+mxlC6IzUmNFNmbbbzB2iIvHTT4GoT
cnQwyAnilVBfV/RXPHGf06/HkUZK+ogOUqWjhjwl8kT30uM4/LQ7ezZkvl50KNxTcYdHMZ2SnpO3
mQaqprBcUM6xva0cj3wMnxiLFBtoc05b1GnLPfzCzE561NV3rcO4lb+RhWGwMIZbdZpNyI9jK27i
ElV97dt+xk1rpB/JGaMl3xfm7Ae21TYVrCJMS1UcBtk9M9M9srjutWxqHXKElBAsRA/7nE2AlMJv
nR/OwetmiOXjQnMr6VOl5poOiZcHSI1w4n6foKSImr5pgUhXafpfEf2I4vtiSMlItgUVQL+RDFa+
8mrB6eIi+F3eP1D2UBX2gc0dcZj4eg6Nki3I7ovsNu6Got6QwSc/SulmjMLXoxz+kdm/Xn98ae6r
M3Bd7jsoE9Si6zHEk0hFx6L8ip1c4aE7ayeVPlo7Q6Ly0wRBEXhx/z/0QhJxms38mHIXH00sEuLp
3QpJJLnaZQY+ZcvK0ZcZ2e2r0YgpSo1hNZ97bDt0bLWJPnZBUEbMpL/PJjKPxK0vSZGHPQvKXkZt
1Ezp5iXwp/WaydCLWC4kD3b8FDL0BNTQaltivM9WZSZvzQa2HZQ+Madj/saDb2MBbjlTsMt90poB
Vs8Li06ZRn7qacFbnEIKODpBEpqwmKRAlPmhQS1uUOWwSuR3emq2vTHlDYVW9I88jQbdNa5ZVeqv
zOCATuWe8Pjho7QlyUc+DfCoicdytMu/1e+ogxNllghgsFCSzhH/aX2w0jRtxduVtXrMciMqpGJg
tJS7qZ7Gjc8xFRE1JbiW7IPo/OFBQLwIOKVH342RuwhSC77aKKOKY3/WUahyrWK6OpL4df2Eo8fK
4FCfAN1AzZw/k7ChacprUlTXhjEdDm99RCiPGLasAWLGleljvA7cSt1DZNHtkdoLjFiv6AhMspOu
NttutPXxL9+E79+CkPEErphRy+0WMIuJSxApKwtZkJumH6JaIF9iH/qeWZxqGsiecCZ3P79vw9Fr
+ZMws4OKwj2taO2HWxH3o6GELiO7DOzaa+/6QxuGiI2lnBN5GOV1/qy7PQSUfGDieUnxoGrKlrCy
Zmqc5g1vRXljcPHOlXT4KWB+GPlh2U9HAQNkxjsLfNZkV6qfe5+Fnxqj04X3SqG4VeYwc/Pm/kZJ
7IDPa6/OH6KuY1mCllzUmftfhSFbtD+y/KdV5IWSYR4iv+BPI1n2O2r4JkE0SSQrlthZuR6Rk4u1
BIMFqLMnlJrzFKhdMizBopOPgKZGKM8yw4b/S6H845vmGYZih3v5a3dZZf/PHSY1G+RgeWfcWV2X
v59Jj8BjfGXMqv62uTHBULbMok0aOzejF/qkI2MghGLiFs6ZigtCAwj/p59oeQolfn+oKjZT0vgm
hKJHxtJ9kMtjMI9Wew3RawjQLUfkN8YBBf2qWKIDpdLjBH18U7fUKMwwMX5ZSVqVi+QQs8L8NmPx
6tlzq+9MP2zfWTa3czNwfOmgQRbZZ7BIsXAwsKPKK4ckggBBWBL/ieTPslXQKXlZVDylCkKRK67+
hPp4EyND+UFXtyUFLUE2uDzp2ncPwvVOdyw9TN5C3RjDzbNgIKjd9jqJtbm4VNJ9Tuq9IYFhCGRe
c9yZGAQ9EcuV+apXCsHXMuELgNW4jmJ6cJAGwvgt/NY/qHVH/wYsiD4zmqjtn9iGfZXJ3bRSVOrT
4520Ilx9cULpMxagFtVbeKL+jAJrwQVVsaQuqsUMij41aJME9Rwiq3s+2xdNUrzDMie6+wTuYg4Y
aNCAs3cyPv2iQiYy/3hr9fisjlBylmKp9SwWSRXLPifUocalyTCnSKTAZK5pa5XwoiTKzltQ6xkW
xe2CulG6IuPDF76SVeMaMQu2kVPf+s7aoHvcHizNazdy4+XoBWg9Mq139/cZR0eXVEhWoVfrYdYn
azf3+9P8cceQwKoscWCsy1es6iR3wXrfknNRBokaSWu66JctnS1Y1ONSt9WIt3mnYOt6zPVcvNnW
hwygGdLSeuivHnWMFfEpCEz32SXFXfd+m4rLbYzoYMQMomxwKh8jmAcM7x1KlQjTuFrLX3A9n6VF
+JhJyEUhjeTJWM4w7qW4IywD8cMxIkXi4BMTPIATkRwz4eGDdFWoX0eZS7rI2mkPo+65td8z2yWD
Zi1wFw/RNSQhOw1v09XEHMRMlc92Bad36iphu5AuDVgEepHDfmSw3qpH0IK1HiQ1WZkiXmkOtkWW
zEU03GXbfbLTE2PMd7Ur85lRiFhnkiVgMNI/JiecYCKuijtA/8lhFnfoSUHC7qiR+NXf/wjO095t
Wh2rfNgZJHn4oaJKO5SFvXnwCgeAXIIJwpQLjWH3rDFeobGEIN0UVn2Cuy/7pnc450Jd82Jfs91i
FMddjdjFkm6QkONZ/3WAbbw65Be+6w+bgUhy0bqQPMwa/LSQyFMcMrAHzgUKdQnkCi7z92xx+35r
Lx+871qCEVQoIL+HxQnSf/hJr49FK7MIiMCn/u/Pzg8UqJSpUp/0H9xfokLAqZJWB8Ou4Akh6jZD
C/ife9Cgj96xvMbVPPSactQdI+3x8hFuuqo+gsNe12RCapcdyPTRColvmO1QHq9X4GE6X36k8pES
Z788f5ohjpriz9lO8RiEN2bU3PtjKYJTlxZCnX1FcPz0bvb4YosPXhMUrl4AvjcpHIjqWKuYBoTd
LhIeGOmdEii60AnT0z/C7a0yNt/q7H1XM9jd8EsjSlnkd1ZrHzmrNptFPmDuva1nrJqrLheETmiC
wJurbTcys2fsrEm+uR8B/XLuAbrBsDpPc0Pkw7R0gMwiu5acOsRm5+xEswJpWm/ftFvVfua8eHC6
orEHhAxIEp5kSA1AuDRDuru+ttsOdjDsMOSG6fIBD/gcw4JYvsdaM6GwPQ02WTqtznIcaGL6WrBg
qNX7SoYjV3cAbIZA+Q5q4sRsM+AsgY4ureGYrmugVuBPwTaRpm9JeI7J4pNyg2bWuGvklzse+wYo
l3IObNdJ2XFEozOK/w1PaT8+ldxpt4CoWJFjrQgb1/Bd0pYvbSYI4ZE9iFPWf53baaQCwh0eaXJW
yxkQ2w+0Bs0Yj3qUzDA7wsuGG5dVLMrVOsm47i/M7Rks86vyKmrbVT+6YrWQHJigfyto61HTB0yf
ULi7WQgrTveEb8I3qURbH3Fw7E/jwQUbjcYfuqY2Pjr9Q6891E0Dzl+ESpPDw6qt1pv/Iub67aT1
0BPAjK4c/QclvlE9B8/ybIqYWjI7Iln8qBMxFGCt0LWg4BhWWoGuWHAT1mvHGy84xR9u16GYQsCx
/kgiDy+5ysBiy7MH1JB608ARolMaSoX9p3pTeOB+yOnbo4RJQUnmYZ/1ZWRzHaQxehRsXwPaiFsG
GH0hzs0+bWCBJv4Id0r7aqHqqAX3cF7dpgwDopCbwrT3vm3JvaPrpkj2vFZkslPP8q3ikmpCv9lx
Ri1S9eVo8EHLeUlkB6xc/X+TNFIC4I+mZvqwaNyXFkY9cFVS8V/xUgxtsS/gZ+Qa55nHwua89zcp
vnOubY+eP7QHKKofSKGDgtUXDqWqpnI8XVI3kr+G+LHzCB9oDExXYygcH+ZUri5t3kV+hRnP7yq7
LkUwlt2QFnb89W76hwI2aI37Aa2D3wev3CRBn6q0vVdWuyYyntct1U/jzceXMDlvl4iLua+tV8t8
j7o9p5Sh8o4zk4GDtrKlpt4RS8VbSEPkoyZIohusPFK5S7Vh7VelSt8DUW0HFRp4Xu+wioSTm6/0
HWgjz0xlEx9ocnYfyye2YHjf0UGkrSLZOs+EDegl0NSHph0JoXZf/W4jRgEmLFBsrHifT6QYvAn3
FOVHcQDBPfPG+ImIrvG1K6AgHDvtK1UushTTMJKlp9BhmDzQkFM5uXHqFIHgRE9qhiODkevKkudH
F7KkHcnQGYIoXUUPGr6FSPGKXJI2EKpzQ5SK3YmLS9YTIwTcpDat8h0WYFHJuTG/+dD++D5t4GLz
nrZbic2HKfjZRRBFIKmmLQXIS7WA8cPcRiKltz21VykJbmH13u+90vrYazkYdsJKOx1E1RI4lPm0
6DhHgTiJqiPSm1gwqD/mk1rq49mJKeIPUnyjhAAW7Xe+la1/tV3NzYmlmbsbT6LC8zr/msfu/CtE
2yU2nk9H666dqehxHGsuRk6GyHiwJWuUdl2mWb/pvFZ8AZNhrDswilk5FBH/+Jb5qwZk1dQrQfPv
PjJSDRgbKWmRLa+2a5Kbc3fpVf5HcxCJy1gzzxR9sbdBZKjD3tnIatIAIGdeaagrrBBuy1e2MvbA
xeJ6um3RcCIVxurUaJzY/O3Dmk/5gyKovtwYfnJKSEkgAH6LMUsUlkkxkCshLTGBv0DNtCz+MoLW
UkzH592oZdE82c8lnAOWuuLsY9/OhxAVWy2Uyn0sjMnR+bMqFmvAEFU9UD8N1kswtkZiUPaVEhHV
Xwy60gBQ3bIow+8lFbIJaVq8/istxvioAZ0Mj9Sri2NrVUZ4gocNxDYwbneF1WkqZJ0W2Q6ajX5p
CXeepm9U7IPAKau1UQZVDfpJH7WSWoezlSwqUr7qdtzw/Dg4fBqgfLlcbXEu1B3t4SIo8siagTjA
6hlDBJ/V7F5WiQfs2+S+yqeZctymTl1o9NvEAE991i/WFXf8NrsZ1b/7UIcRzt7bPal67hp+Sfha
CuuiyesdwEniYAFGLvBXi98KpJl6ojh03dhcQs7wbtGyReb5vOqGWBArXdYy/EnrmbBLOirnI2xP
5bYaD4I/wpRkEeTfn3wAFNzuNht6PNqsiG03gp0seQ+5trcQa04bzPPabgax6u/eCyndbFqPC/Wd
JcDVXGtc01YcOhYz+9WqK671zPT3POnveQZwqrP+2RCBGtYDE2GbaHPp1iv7oRC/eIeLI+CEm2Z0
JCEg5gghZglXH+5wSWGXornHUMWuBj7GQ3ng/lHEgQhgNfTwfbZnBuMJ1LTs1eMpawNOhbBPRF4P
YjQiux8MnJFtZ/tY3GKC2gTUzUZi+E9CDKDl1QKkuoT+YLjKdMfVw7C/GVjd9Jqa8eRP2P1/Lcu0
AKDo3Uk/k0G+Gxeno45wVMF2YxASwtfeU9oHmC8xOGsSQCiawMnf4fEwZk2uxpUEYnZztHc6Zhaa
aQ/4dPtxfnctN4CzbPrznaflbgXBs9JeUjTROryDt54/ORNZNKK3/zKPUnIIksJJg2Li+s0BSNJf
5ZduV8f1WDzSJ9LFQDEUv4L/3VBSVGRhRWvSWdiWOOFYQLZknAnbnb5v8/IaSUmHcoi3tKOHXfS+
sIgzr1f6S+/zKewtDBgUWMidAiE3cn6H1ZzEP1BqebQnFegexzaEOg1bWI9RD5up7H9D1m75mhc1
Bse/mjzf3MFa65SICdea2ACV0eX3IsKKHqny6ZfrXPnlfo1YePu7FkxiZkL6p6gOzYkTNfPLv16/
X44ReORiOPk7xV66si+R2tVLx49pjlqNsMgX89C8Ke8WR8EzYmq6+ABN5TCqT6i/Xu24k4ioJ2cf
afdn4WIV9nN7xlAxHDwpV1X6j/FQ59OBDr3Y5G1RL6SWK1LfUcvBV22GqCF7XIKxolAUEbeHSVqN
9Ps6pbTeXd+XJLoWNiwASrQ0AiS4OF5ohWPS1rJArnitcyUylgGcnQw+kkRskANLlBL7pTtkCT0n
mVU50a1ZKjWCRmTzqQUHBf1i+Ekg7/Xais6iClo3fGlmGcBauivn8EyN0M1yQr9pNJcnf+7F7aHM
ZRvOvmwICtPNskDD9LRxX9/WQH4y/Z+ZcrfbX79j0b2JzSe2t1aCUXGh6dEppZAMUjEd6IR7f8uV
VMtfjKZFSCa0CDnWERCfFs0xg69Aa6fQTrZYqmtY0DaeV86HS6CADMQSaaV4k5wjs9709ED0DpY4
xeIzhHmHkx91nIpl84zrkdcR2a48vlhMO3EA9eOf0GLYVAKjJyiyIDNVoiVK7ulSx7873wtNmtwC
jwQ3d/4LuWDVXmK8+8XLHeFQMTQykZccjWMpTRzB1Mg+JzyF2c4EecoR9SylD4bI2ORnYKl9Sb+v
YBKkQYPgz3wLdPmvjKf3XEoNny+4KgvxYHIurPky7GDoUjezy3XyH0nfovRQOlDp0CsUk8sEfBxc
pJTv/ntdPVzB099fEGAsMWIjJJPQYQ/uPdZhnyN6cF2kLpVN2bj4ZylgjgWrDPk8zIN1EFhb6KYN
g9dSYDXfe24wk0mWgxKns24TCUbZTthBouUwryzO8DivN9ovlFBgb3eWUAUweoZqLVa2Mdisf+Lw
748IUW8lE3SxkailjJjsx4YxkVlloRBpJUaT4IOd9jGI2AFVqvCljE5FSPgzTPslEy7KlsIaJVA+
g2YdvPmEhyYFcxEnF3/adRxPv4mnLrPqsX0GvmQqxIrsdiaB/qtQWv95diAvqxxY/xmdF6l+KTQu
vw1USG61+Tl+qwlXN0TxFSzggd6oTXbRsb9CGJgIjRbCJ1aIq/35GUffNCH6+dollXpnvsgVoV5f
8uoM088i+QXewgmCyY1hDwY8SsJnM08e4wVNPaJnc/TLJC1WLitebOjV/sNiqX/E/Bqjt3lqhbGA
MP6ubMVeSyZ9iG/BWyYhVnmlhfB1MyN5elyKMRan/m+Kv5V9elboXTy7lsPtCE35pd2qKiTBd562
DeqyM7aZW/Z/bejw0k9pZhNLtLVyvfoJ0G5HRnqRYaHhhuYyaYg9xdZdgilpgXDtA9DT2iGR5FCF
T+C9AlB1YULdMaegJvkJjDB+Qh0y9XesdpMB6wRjw7jnnRbACSCy8gkwdXuYE6yGNd/lCU98m+GV
58gR3tIySQKZ/sbFGZtt61MQnv4skg9AQ7D1c2/wg5ODV3GCQifgo42/b7gxJXftn6ZTWQtUqJ8K
24ve1VkGR20MI7yRgJSSCOCK5CqTxwWleiMmL9N3esKEw3PkHGX9zVQ+TWnPREdIJfP0RWE43AyI
XQwUf4nmloa+TqefvApxpBdIi1i2gQfudtRG/4X08ggumGZxT/upQNy2/rP2zzLAihl22ZyvEtNs
DuKqy6wBDNO2oq2ZF/o8HgIfP/E2yVxYpV9rxBdMteMKcScM4RiqvUMCt5eOENMexKEKNEclAT1s
TOhIep9TklDIsKwaYYbX7hOt516uaCk63agslaG1bW6MPqw0ZMRmBZT3tXuIV1yIBrQ5wLhGqxL8
cHnCdcxYFmkRvfrREMQamqrMBBS2tT8MILfILGnWwdhG+7pxD0f24h7XZ/OpClkp1UOtqsF15ZWO
RYxrENIXQJGHwVdxmf/Gex0PaUNpnIm4nKTsdeNT/WV3NUfkEwUNOQI42/HmAGFAidmbVH15IymH
WT86izuQV0kcwYczf7ApLYzFWVaPvdQngerA4Wvb/iGmvWnCaQq+T6SlpbjIHU+MIS4y2ZZSXa0z
fftBW+3l8kdLOgYCuj0JDKhJOiKuZBfmdfsIHe6eLUlrnwdYwDYAswFMOP5JW8bhVBuEMsDJ9tvl
IEMDt4CplR/6A1d2hzBqago5Z377CuwSjuHxsn63v3MmDuvqc7q9rcXJcWBD7bl19Swi2BvOx8SN
sOsCWVdlxz8oU/2WLguxWzXHHkRCYLW/8HdPW13Yp0FZx1KVqlYlt+BKjqH5iZDV8vfhKz+TW1ux
nKOuJNSCq1/aZ1xHzYBwI/djJ5NRBdov6hj0chsVCBYzwkJOpwtXLhwKIc6/qvjszYI/9wDJjRKj
0008lKQgaSJKgTVIIKkY+QaiggYdKLNgbmjRGKUObswS7QJlK86XbTFeGlWSZk3Q47ik8jtuHS7y
zADcSEkWHpBwTJvhP3mRyFSrtGZdRlNRyaa8LNTi2uqDp1uV+gJvkak0TyH0YOflg1Uv93FO4oBc
VHgHUXG0ykZTpwSZnxuoCIHYneVoXt1N1vLdlcCnfHmFcJLWzy9ytLvyumIDS/lHFb3Jf9qfCmKg
wzMoN7bUh263B3SJnqmAlZaW5DC6nw0rbEFII5BCVwFUu42XOgdRG1FwlWsUl25xDuEFxm+GIysx
j5ecAkEJu1EPuJk8pQsAs+ZS4LLLs0A1NzQQDjz/8K74oq17zb6FDW2vs/lpBgbxx4MVtHIhJ4/S
phLc8t26KabCTRy6WrwQtSPU7gX2YpRnM3gnItIe8rflvzEVQWIsk5iHhWUZ4xB1OEPBhr+aU2ju
aQErMACSpfY4mVECrn3R2519HRLCI3Zsv5r5snrMTWrHvnnYwqVogMZT4lDI2h16uVl7iYmEngjY
ADpEshzjQfToeuwXkX+pdM8KyF/0C6QfOHrJ7xXYRhWQ02Qk51KxDHybK9yco8spz6+i1Dr9YlUz
2SJnzDnnHCeNjFwcKwrUGLAcP8kdHvymei7U2GoSfCbnRrdanE/NRASpnGmoNB/dFlpluVoVhB0h
4i23pNhFmjzZp+LqRvkt4RPfsKmku8wxT/UVPu7wiL7KhlYIZvLGCI8FcDJ+rRyj0i06g+fH+96w
QUVVcRL4MS4ZRhi4NN67odAJTVJcnrPh0rhEYwWcH+3YYzgcFHzYkBXYC+qt/BwBSuUltm2FnVRy
iXY99TBU7pwhA2pgfsTy2iD2+6HDdcLbALjijp35mO6JkhU89euseJpWCYbBmkFjC96P/KBS2lWP
8lJOxozhcaI6ELRRzIdKQzW1JVsqR/BsgqeW5DQM4+ErKttmZa0aogWbiG8lDb3WafY17CXoEk3D
TdeA21FjPVXEZaB2Y7sucPIuL9PGUDAFt1YPdY0iRjqVoOry+QuqAjHcZDzjZc/rStRMYOHh/lcc
MGGhmCb6pO8R3iKTYiluvOAHJ/7+rOAwKEauD5dHjmop+8lWe/AEIrbKIA7TAQyPMmw6XLmfgeI7
A9r4TjyYy4/cgIeloAdL6OhpcWsnEz4FKySRBNyhWmOUe7KmB/QJQS8EhIQEvtKXg7+TTySxfxMi
ntst/T+FB6Z+9MS6xXySMXJ5FNPs5irtUXYfb5wnUGTxobf+lD3W/P4i22v4A20FUfjOtzm9eU6A
wr2ZFE2OlaLxIXxNV4IFDleiSh3Lqv67DLXxw6XPpVvG9GL2ZdK5rQHWrWXVdR4D/GPbhtC0efoo
BjqsJ4JVdxy9czIoqDloCyVfv5EDnTAtEVCeOY5GD8R/nG6v2QivqTfVrfBes5Os8INyLYZcCiVN
px8DsJJYe6hnhWdxFo+0uBIDfnGm3jtVvLnJdzVETRol+MSGPwpVo1xHNZzJ+Irfk8JYcUzJenGa
CGYKp3C7PNgFgFlbz2XOGnMQr+ASCTwOhnc9Y/nS78BoyTibpe8Wp7rMV/Q1K1QGlc5hBaRqdnKL
OBEHO313IuMDCu1Y0R8Zg+hG46ZyODCOmCzuLDjuZ20xdRyW8JaAm081jmSafr4BsqTJUjUa4MUF
441fz6pTu+P5LMqYi9xbUzbI/LvY7cLdOVqKWyjE7y4/X8Sala05Z1f7TzCZ2prN9+1YF8aEWk9C
Y7nUyYVvNMYFv2H7q2UBorw2UqtVS4HDhwfzavm1jz/zr48yNTI20ZIfQKamGJanLZ4JEw3U29cK
TS/DRsz8s0pdBbPLJDPoHN0BaqC85CBmjcNOU6hZKypr1BwP11NOPcZ6zzL3slVSme4a2CFQRfGg
bbCwg3NCRDTObddwD7NmH7iYvRTYetHCftjuP436HNrf+e7QHt8YOBj+ASzRgF+UfBUzNPBCR2OR
XH4oyuBJ94voEDTyzfHcI5R7xN9Kv/hudo11Z7Z7jbwGgrHJ51tC4tt/ie/QkPGzs9pODXuTwZoM
AFDtHKVXLtY3wtxmjPVaEYrUsIxNfB3qIFtTluaKjQCUxvqjbJzx2khOaeTpAEDsreNjAN5E8kZF
TREnqRLtZ2wE1etTHrQpzAKXbDMyqvTR91taIPc/lm1rFnCRLCguNfP1aUdcy0YL/eZKNWICzGK9
8X/+Qw+w7CRqCO24XFQz3IasidaoEllHd0pzbQYZJThKYs17DYysXeLdKdQkvTwN8LuPgnBrHd+I
8XmZ6OaCe0ApoeN5be5jDSXLuDdaz5Xbeq3dTQNwKlorwCGWcSv7dXvVGOt664E2YetpcLzsAELc
UgqD35lZifTYndy/opPG6lWuz5r/E7RY7RgVPvYAvuRAHRWIjkz9ODRMDzhzew8ookgjhuwn91JT
eFatu0QvqWP9JyiGMuluvt2Ql48I/Aqhv8bbh9r6oU73kdpSXfmEbCjeRgTk2FAY+bSDZ+14cu1U
ixPM5EaNeBpF623QL7GWTry19Rljo+yfLVkBRESgkgavaerYEUgJvAY4UFek482mxz37JFpBgNc0
0j1AYAem5DgnfUsKxlyWOj46idylqv1CezRKGk1k4Cp60/uefrLtpiAEAgvAFB6QUfV3jIPVd90S
yobXxRXhXcifoLlFMTylQjYKAtUQT/QEyyqJNckp6xeXgi04VS3m8RlDUu7l5nXUqMxKGVPhF/h9
vMfCWvx7HD3YLSro8wlgPd8tWLXLfEJOQ8apgcVSRGZ1FPcqT4L7iHKvXSlsjsyPOFM3zEng8570
9b3Q9N/Vgs7T4h7PXvVErkgvmzeTev57eOSgWLmP3v+OGYB84bKKp/x4X5fkCXYSGV779RxlqJha
NYQNR8a/rAKavrohpJsukIcDnxC9Z1iKHvy5cP8KjGm4+asAjzAU7ODZCQtTwBCLMaLmceyZTd93
gxocAMQBl8G6dRVG+K+/gs5m0K40BV9t99qzoEC29Eh6XJSBaGlcBk+2sjOpKFHbJcFYF3Bpxesb
ng25+CDcjk1QGhlKpUm25tjtRugLqF/NUMPSfYfBjBLp/k05OQWuuqRLlZZB7gIP0iSGBvAl+eX5
rx1O6Ay6XSMyxTaeArqx6EWoTpIXza6SRuR5dmxHfsWyOmKUqcS3JTa8rZZJiJZk/HO4jtL/UiGM
w51jfAd+VyM+cEiMo3O2/A0gWS79w0LS7x7+aOcV1mh9grx3iV8z89ntLZ9wFGuxB5v7Mp6QMqfV
CXAIhkLitKCPTyCY/MXoftNOnEA+jJAxzGE7heyZKPCwhP23n6oF8mm4FdOGBVrDpkWFzzKDiOBp
SfgLfRYL4CQEqpx4VnghyUjGaNmZYFiaW4rrqzEx52HlJIgLON+WZLx26kViu7vgWhS2VST5bjy/
ok3ec6IDTV8NBUr5IGLpV/0gtjJSXvPj4iPJcwQ6cRs5AqnfnQlcC4TePjPnTU+d2Ucut2yMIqIP
AYZWQwrVjlBWp9HQgFahBKSWKw0yw6dG//RSnPOUABh3PomifmsxE84FRRpqNVn7UdSLisulOr/g
M272QifUupIGK8707RQrESLU7ib04+7AqVwtOjcUsDm0oAJHqqhJeaCCQaLs9hFiDrFWQtO4Jukt
97PmisSKX/BEsB9MTXloo4yo5u+T765SAi/49NvXM9HvEDFL0SKl6pRp8BDJ6TSM9Mi9OaEOVguo
sp0HSyXLxK9RKWonsz8cesBBg0MM3yVdNVySnM7PzxDQ7UWQaReG4+jswH32XWd4hPC4z57af1mi
gebFPwug6S5I2soAXgF9Bw5oYauprluabC0JZ6xZYskDbcXOQL3ak6dJ26LrvxRXHtnHAbOM+tk3
RpYmrmuAsOIIqUas7uKHXhbFFBirBMBv3tX8IiBbYjeJD8KFiolTCly71F3ibvJCX+VUlPJ3YncX
8HNtAYioExQqM3mazCLTtwBAmvhVN6sLoJt1jUlyOTIlPrrQLAs1xf3Zb/Incf81RfvFCjszf2qR
NwVZ0rhyp8zI0N5nOufL3u/KBCxYtUfWpRr3v7GuUxIabxiKkaVCDzKNl6wd51YeaHZsQm4JdynO
CTKQ7BBdumks3SqS4QX1T535QEsPbkpMGmP3I+2lVoWAaF9NK6FlyzHpzsE7apoW663yX+CBRLIQ
eGcuQu7cxrLoNFHZZtgBU0aRQ2MRff32w2RkkOTvfl/XhKEqX2vz6GOdZAX0qS5zoyiLw2BxefHO
tJxutQ3Y2lUykuIrNjjcBozHMKXvRz5yHl0FIVh38qPBpSCD26/4Tnk71UGVvGrz2fX22jfSeJal
X75D4MhEkRy+abajrcxILkkNfNlNDMzCQ+JosmxIrFkWy5xepgFe/RgR8IwZ8Evn9yEuZ/zIl0ko
5wAtDDv3reFB7vx5xDdDfWz089j670A/OBFFmxephrL1udQXTaE+kQZnNH/mWHQYddQNlNoWXPi4
WPGYNrS/J3OHFyQ2idEUv3BEUxM7dF/Dm/LlGLsmpDAn40A0hpaoDI221XiksyAld/ddN3vuwNE4
Uu5CXv1p7ctxmmXqJFUYaqNf7hU/EMVz88JAP/fUH9I4/cCEUtFyAbNCa3H/6F1xV/YD649O/MkG
HCcotgDd9dq5h6+Dmp7S50hskl/nefF9t/kMzql167ipUxyuJRFm7k92uY3xOAHcnRLSRm2GPWh6
sxkwdxwFL7ZCPjrpeqf094WOSqbpz6VLtSMa1hwTz5/A34gcogWVtNw7OOchHRRZZBYbT7QvRM0k
h9G84FeCL1dym5eLdvyj1w5TBjc53/ytMOn3uXEVFKzrRrkTGfgrOa5kdOX/YAfoFlkhTy0qBsEl
GLX2ufJCvC8pjIjJiqPzV8GrrRVJNVxqEffkTgu00fCfEZ7G/dv2K9XLKBkxENlxIWf+Zej3ebYe
1c3tNwCqKvUEVHhzqKM5nMVazLVb425gAX+XBeiUr8C5m7dZtKq9Pn49ql27KHJYm4NX08HpfYO6
ylIEICJM/lucZ8t0xvUfL1uqIVLPv/GUBU0+uHx7E5XoausuVvSgU+zuSfvHF5jj49i+ZVzH7wxJ
2GrkBQDdIqO/YUwe4NloVojDFSFhY/F810qo9YLVPa5rLxJF9krDk3xHYv+1/LfzQ5OMzVh5R46n
tfd1S1MEUcpx2INBIW05OAypyIUz4zZF52bveouMdH9X0BrQ7JVf2g7BWl4cBDpm4p2RIj/ZCb2a
qvU4L5xsb5K/5C7/5knYj1uHXfnr9ZmNaavf8MPwK8C+3mQsczJjfW3ZE+dZNXTGDHs0f373qIIn
L6Rp5GGTpluMUvHxN1AILfHGN0ARtwt3OdfDYS17KQ0mzDn/5X0MC+nEfuUP48RpMWrGz0QLdznX
FcmY3HPRC8DqZomE9c9JNnb7qXogahocKgz1NePnu/+rPMIpP8sta6HMkEHirESz2aaKnkZPTTIe
j7MgyNP6/hb16U/SDN3ovVfqcBX8ZAeLbSnmcFPiQtBxqT6HZejbEgpcrovhiLbzRKlg4BOdO+Q9
9RD847gcLTpV44yFBX3NyG//XRF5PhvUiGMCRZvRR+v3y022/xUv81acV1FNbkopuVcr/KQud29L
yx0vmZab6/VgG2ljlYxl9l/LQWD6YtUZbEq4IqJNKwUWpBYOAzcS4T6Qh1rwyDUqecCp15SLGDI2
U+H2MdyJ4S4fOfB7lrkQBz8VZMl4aJKWAJUqknLRxthG7lA1Q6ecyYqPrBkOOZ/xadOU/hM8s/2q
RCEBs3WpPyYh6uv2OD9SHga7R1OrDKxtLRsPo2VtRq5VdkpUUwZC9dGWwxbsooWYjC36Oilz+T2t
LtMZr1bhI70IXTAn3ZTKS+DjyMqyvd86eBMlBckxTqMbyDlZw0MzB5D/dVVJtM8qEa5xHrEV0Xj/
1bvxL+Jee7G2R8aXtvklyV4wkf/mNxyrls57A7ONjN9ZUvBi/8xp0QTeI+9s2kUL/VVElqKSDS+5
WQks5tb1ic1yu8l0mPKaaozJ72XtMwtja9km5+U6Nhvf/Sk4sIaSbhHSNtGMZRD9PLzeEKhtoNTr
2rt6p+Zh+HWDUGjWaXce7Py3bL39LtBg45I6kcp3vtnYwrxGCbnl4eyi0Gyr+pEZnNCUJFDmNbny
hxTto5nqQLAwAQGdnBDbem/5Bn9BqagWM4iNL4ElINyTiP1HRYNUDP6H3oZGEdZDb6zrcFA+JYfd
klhi3LQv1bSdKz6O+VxwF3cwLbWchebUcY6tKda+F/MqQTnTX4TBzYS6vH6sVssfmT8pUfgE0/iu
VEiwg0mjIuEh+aX7Ss6kPE5+5NJbwoeSeZvIVoaacaQMfdhSwiWWXzv9wAQupYH2nCKaEbsQi5IM
BJ3fOJCcRYvTy8R4uNjcLcpOIl9HqH6HnjMNwHkzZz/rZk/r0SlqEfmIFn2UceAlAkjtZkmFv4xw
y00m/k+IFGb897fRAshslCdvRUFe8m+NcBmnlWMC6i3X0olkLopsJ0N2/wEKWGYCjVbzkBSb0bq8
SEallphMM6lOWXWe6dVsa7NroVktc/SYow0t3Ruu+MdZRmv709hcWHbhMpO6spHi79IIPazmKj6S
kgVfgEyUj2MmOJiECdtuKgFbciLRmIMDZ+h1Twz1OmHyZE27r6pMmq75JTaxfV19hkd+REuyBS1/
PuHxIcySOo3Hl4F2tikU8wVlePkcXe1MphYn+PJ6nc5kkT4FQ0UkPXs26geCjKZ4J1Z2MJ+1Wvot
VDefX+0/BY1+ek6kV0ZAmpBrYWZ1U34NJ7qWF2yZm+QWCsaSXotKcCHrJp49bxmv7SqijMx2EerD
KNK6pToETQet5YcIshiFf//HdTm/C1/Jiea9HAsD9k9/yzoZEQxGfENEyuoIaxBU4xWbfwd3MC5T
X2g0CMR9H3hFjekbXG46FoHID6TP9tcrzeWUO/Ngd21fMh9K6HFOB2pVknQAUgpkMj/klb1qplD2
IvW6Prnx+pvfJ2uTKclRc9Eo0nI6uXMHmRkIRf84Gu4RVsTiBYHzqBXUjcKYiFDQSwZKtQQp4L02
iFVZ1ewE/O+lIVX6cKYFs8kEOq52SKJKSCTvHyOgVf/BsM4TJlKol6f94QnrD6sldRW5+rbVxxQP
9Aa0bbpj8AoliPqE5sHwn501OwbtrSws6MJx6x6KdgJ0agDFxQ7Ag78WNcGiR0WAUgy+3Bw8UglO
FjyYm+Ko/1EMK7ovOYp/kmLZ1kk91pW5WpCBVJMKBE4LAOLXHKm2uOK0WMdBeebn2ur4C3/mDc1W
PTk1/b/8mKngdCoUi5Ah3NdE5YzrNsRmsxqoWN7Laa0UdXT76aLdjnD24GZN4ICR4OnoUJTCEFlH
QjOPjbLtIjo92ugt5UwVjAiog5tu4IJdCXrt9H6WoAJEcOBlUvzgTV1Lg3USXbdp3OwTOzM8PCa2
D6jcRgmajdVzPs0gHehu0mCcjjyuoL6OtWnlNl13SeueqBYZBY0/2RcFilbhRDLinvI0p+GbAZfy
OIJDA0tFL5PxpChsY5g+rURhFHCkCcHCCYmNbQjtGBlyYFVnMe/IWRqtQtOlGxGQ78ZMr0oQZ1d2
Zg7sG+Q3kvFYlzYrNHSrIEaFA3N0N5v0peJvDO9XVYSwcUjTCWVZMrDcIp8q+h/6tem086vvH+VQ
4eLu+ADUMB2oHQ11VZuo2XIJbPOxvSsSiVCaPgfJvy5gdTwoo9dXPgmOCDSdqwYCfVFg7qCM0U97
mrMpE+WY9euFnCyarNEEdR0cogikgHQzZp6BVQiWj8mmI80agQhINC3Cq6OO/jsOtpb2aiunAhaT
JeCADeNkhVAdzE9XeIyvt0oB+q03DR7j7ocqCTgTv4iBjFzCbXQP0rtu6Fy4gF5F0Q+HdqRC/sBx
sRRYA6aN1CRED1DDbN6ErnKQL0oA/iPNsF5VpgzdjzlLrTnDT7S3HPElL3SuB9xYCW/IOYFRjYhn
woX5cuCZJujb9KXwnta28VySQtrIlzWIs58ZJuM/CycG2HCIoQG6ZfHpak1PFCinuPtFX2t8HG8h
3NRM4haN8edcqsoGnPDAp4TC5kNTQ5eajDlOEdSuudBDL4sicrfLuG3zJoxbXFTz2bc/xc/msfG9
UYzbGQBlw8pFH4vjgU3WA/V9VI1qkQP0hwEzZcZaA9ybN5vvsVleBk6KJ1uODZSEr3Grae5Nlk0J
2oSLXVGNtwiuQh175xGL1J8D24LfmFz6hV80paROvkL0BrJPX4C9s6Cx8SXSR1wAQ46hDOhZ9lgp
kBSxpcE0hlqdIVk3cOO9Jm29uKm3Dw0jFSvnqSVhCeEodjA7Z/QGVGus1b/fPZEFCOyGfYTt9AyR
IX807w0Iq1OMu/2oD6PkmdlToqjcIwFSaHYUs40YhqoosLZIE7S7X+72YJ98wW40aegmxBnfezsB
8vGKxxYleQoCewWvgzL9axkoTfiGZftIY7xUX8vwcg4uNlKdPCCtv2HNkgTRmFKW2P9WZ12q1Lcd
KphDc0/O4cN74rqhsGAgyoJjHO3r8p6P5H3wZ6/BoZCBylmd+aaU5yVjF6Vz6xldM7O1l0yK8ICN
ovSZSQ6XdV0eMQSNVJpRh+j5u81JGmqN874CuXGtKLOH/yUpwk2/3Wa/xW6tbqd9WvMA2zMNLHkx
xEmgmjqENNBG544bR9PTI3/Q2LTyUfgvxjdzT3sB6Ij0Tbav83GyGv0v6r73YHtFo2mJfENn8twE
e4hQv6bDma6A3ZUkQhWfzbRzlSsOjGTshBWM85tXbuLicAW7Eg+GUhh4HsWzgUPNKwaeemR06vG7
a9s66TEt5Roymgb9ee0aMldctLNpBy5+lJpirEU8/6MLTzSC3CTBlq23n5AsHfB6zztQTUpq+Pi8
n7DrTglFMTbHr4CIpz//F+qqy5u5ThP8KW62OjgjYM/R00YwQ9fkVWMPqNnITdJiJp72PhQrkeV0
qc28MjcT25LOJMO4Aeq4rZJJcRbkl/msINjFBbG/UkxN7R5Mc2Agdfprf7d4ID4nY6Fi1wufQ0h6
nqNviU3qvbIuuCTQmsBnRnxrv20Z4+Xy50gbqAm2578J3or0TGlUYlUc3tXLIZHZHLj8goibqlu4
trY2Wd5L83kheOi5RAt36lc5Phaxv213DhZ32B3hXrk6tlBkN0WW/0lwnQhZ/j6GYTR672VqHfE6
LdVTKwA7wxSP7u0z8vCL2JJ0Me8t8CvZEf/TjfFX2ML7XaU0owKlrG1F3u4dM8dN0ARwjyhbrGhc
XFaZRTTqgDUpGiuxQ3PTxvv+PEGHvA02DBhadMO+kTKjSERBGFNEBiRWa67V8jseiyjpN+mXS4wm
LAB7cRpzDBVT5f2d3pucA+lgNkh4Uftgtcpw0Pp+K4zud/3n5EC7bqvPu9mOmDHcjHtu6oc3qD1B
OxuAR7pIM1i27NF61Nb+0G+8kJx69mdWoky6/MwYkSP33AvdHekQP/LimtnwJCLH0npBba+/7rD1
XSsfFeCQLKA9qT59BO0IGnRLMA8qop0mxOAGF440AQqqaXu/3G706lhZlD7GPNeZKZmnCfhGyFjW
x9Yc9TboFIJo5oSgpxmAObtPLyFXLFvPAdij8uvSw29MZaypX/i7JRuB+GVsDJkT83Z0A1wWmCCj
8gmYIO6yNF5lY4TM13J5fTNPtSTg+XUeBW3wTT/HY1X4OH7uXYypD/ln/oGFeE5jJ0HW2QWoQ4DS
dKMIumMLqHKG7nx1J4bZX2DxP8HRnRkPxW0E/6eOFLwN/8dhXsoNRepYahBifuNpLUxo7Zt38YVD
bQgURpvzNeOcfRNVoRjnwiuHzXEILEnktMLHE+shBKA4wKDno+H4KawavVpsEh7rqmmJsi/YXkdt
SHUwOnbxuT3oXnHytWE/TiAmbEBC3gnpvr27jKLGmikPrLYnswsilnOx0Gsjy8ikPgjByTUrSZ7k
1vRnABXHnPaWmHXblitd3MZj2wDjhb60p7qWeFuRXMCf5/lALsu5PERLZhfyV6XCpcLTjRinOYcD
YmXMkvo+6uerCUppg3iSP+c9U2j4odZE08TfcLtnN+dHnUnG5j28h5MMjQpTE7TgittXj7ZjhcIY
h3LWKaZSbgtVKjOmckdQ2xh+ak6nYrl/CRgqOA1eEy1DAFjme1lKIMPkDwUMJrRD1BBRnc902STH
8IbL3FyUslle6PuMSBcQaQgR3du1qt0b4kb4miLMtOpvwzoMpE1TVljg3wZVzA8SCXggMccDGL0B
mdPhsyJ9TFBX+P455fwGsnaapH1Qs5vogWVS9k55y3u7ILf1GcbgfyMK/0XpyW8J9TyFZUxg2QjB
lW304wRoFoc9Czea3p0BP8QtpTn0hFEj4e3CkPe2D2foLbeim183SwYZlt3Qt0vfcI2btZUREH/b
Q0nUIo8bxWYkIlNyg8qXoRheXwlgW8Cp9laCysSczWbLsxq8ReMTm0RYoswyfGXGFFg7U6EtIsTc
loa8tlsLktFTEJT8vnkUsh6XgKuDEkxvfMWY3/0Sqa7SyjmjOR32KHiUjRTJr8nmrAFB6eT+JEq8
zm5hCH3KigegQzkMoy5NEVmN1NuFzHFMQ51z/gvJmsuXjHxc3R/KO7zCd/bOg/dawFNMAP2kO+yZ
1bhGQx9f5cx0jHa/cTp/V0fuKb0xpLpLAwEQdmg8yioqLJoNL2jeHgmRnT3X3Lq7ej972ahUYZra
gP+FtbF4eUAn7oNMZNGZPqQxwJmSaqKbW7dFb/AJiWHQH1EgAwj15u7esJKJcLjpe5u3R3rSj4cd
5OdpR+TMdz5feIc3XRhnGg9ZDKY+y+qEhhJ47/vhNZdV+9AvV6okQdHuoeT6SZTIy/H+93p5KeHC
auGPuJOULNBH9bUkz1o5fVS+d0T/2W+Y+T1upBZUhIXuk5d4VMLh7H6ARlXxvxOvS2ya/EGfXn9H
sSAcJHK320AJJnWzQdAG9zeOipLBbPKBp2MW/WFFMwgBv1iLvQU/et/d0PXVuDdR0v+ajFi0Iq46
yB5GU0oS4f2c1FFKzL9NArvaHaa7NZMiDQJUR6zJ55glJGzt0i/UtU2nYD+kF4z6bumM7bHSnw5I
GUEG9xa4AcWTMsU98hObHlMxpCLcEyfg3fghQHv7AzzAQdF0llf3T/lAQO0DUBL6PvTmH5b9uJrT
FbzLGYlu4QOfAaNSUmjskkrACcWyZKkHCkV9stjn8EFcvStllkBvRF7cMAsl4McYCPLSG+f6l+gW
bykiGz3fbFj98FJdctWoLOdv+SETA8e7j9YLziUMQGkYPrHFQqYwvX7cQ/sHcgX8Isr7LkkRtney
vSA9FHQluFALsZ9l1MBVq7fvEe9H+xY+Np/9EbbNF3fRbMZOZDG18ChMyvQlA82LSa0lQhTp+o4k
n3zwMRhkbWR/6qwasViUz4W7REw3R36aJBndMVRywk+FgK5g1xREePo7/1NLXbAjNeFi4XrXz5DO
aUmnw2ONa9ppYTw4nRKcuny4xCronxbuqCelv8a05s+FXP6O/0zZUJcnhhOMwrENW++YMq9faySu
L/8IpT1lrweBgYfhyrycGHJV4sjQJbXyFqdAipFM3NsLc0lI5DY+mmdXPDnJHaWAIIuxSnmjrpyu
Kv/S3AxgV9fn5ew2jZa7K4QcpXWLcohJShOsNaTnlb/d157+A3c49KzloM0xpGWUZjzNXixPR62O
CI7D9FBv4OfFm9J2HRK8dPai11Kk0rCRdWb+RUgp03j4P7AcTXWeyw7NO49zQJQNnFZgABsC5eFZ
gS0+ajFV0z4hH8wbQRTripyunflwGt+9FafJ1GIqQoipPtKsdHfPKTyqKYbhNYkYX8PpJWZZ8WAL
z/7OVkBokqzmExyjbquEbi5h2XNpZrVnPt8V/YkrW9QqzWKr82fJyL8YWLyblyIgUNIEjnOpUq0y
odoPTUCxf2mPiBMXT61ky8vrCjbPxgMHU6e5Vi09G5mOOoq6EZD13xD6mF1WOIE6L6Yf9dtIRdkG
OUh8eckTeIukvOVRAThJplKdy+M7DkUH9VIgMThmCs1wphcTgjNer3CIVkdu1ogrT/ky0DDx34GS
uAhWsMEHELq1COAATSoxKhkfaIYLSSUXVpz8ZCpFoQ7AqB3KyyMvJ0JYgruFbBqZs7wuqu/gCMuB
lOI9WKNZXpQzd7de8pGJkZ9SBp+F3nsmGgtx41brdrtunQAwGK5a43a/mh1fY2c82obu8h6W0nt/
OQSk5kUS6TsEz2194iNZG/syZ4jFmLCy/G8zsQQKq8bBqS4FUxA26SPvC4LSTznN8dhMEgHo6Hpf
RnqU4dzA6m/M68gd6/toQaYLcQ4/mcsgORBa2Zrg6vbe0awIjAo+hEl6sDg4gExkbzlwcsYw1hCQ
wlo0CxyurCzb/JON2jbXPdMRfd/QE/uxQ1Os+LOGx26XlagnxtHKiH831JIuMX9yj615J2pOVsPY
DU7fXlk2UvKyz442Fb3y3Rp7lGVs+j7lDfYZ3gNdMWOqn4u2D+SfRBuGUeyLPT3na/HbPK6eKITK
tt6C2q6tAbRFAryGVnos8IzyP42xg7dM/IGtjnz2G0vDZ3LIkB8wYqFhdkTpKZjAvKhv1tx4ecE1
ujRVQx8ETdw/Fw70/fF6ykfTE0W+wPl+18iTZP968ebB0Av3maVNjTI//T8G15r5biDsgVYtKS+r
la574BTJ+GVVpVCe423tZUJW154AhzMxGAuuQnmhcdHEv+bFnsscnoAwjcHaKIoCtfESzBcxmuRP
NDy/A67rs7STd5nogcmG0m9k4OOz44wABmZW/2KPzgY6JY9Xq0Jbv1K/NKSZjOuu/Dik3eFcz4GD
BC/bsspS8vwTY8Yrv7+OBtnUu3xUYpjEVJLdQ/o0rX/sGecVIK8R938JxkGllaC8crxXhvyjo0mr
U0rUqpQYdCMq3RbkLpfGuVLQBZFQUI6wMnhSWJUiRqq3hr+yAPtWzQTrKmSj3iy3aN4M/HRk3bvK
jKr/J4RySLOJIewNG2o/915GlgGa4/dpQHNGd2dPnpDW+bgx26gT4kkoWW0mc6IGiRyCrMCzWu3/
ok4K3/4MKnbz74sVcdln9FH9fYXfsIck9inzSmWdXxYd0izYeq4f4brsFYTar/qjo2nNt08h+jGi
JEY9IZj6Gnt7VJvsEEtxIJv0bUqdmiTULmd7pbjyprtC0vkNtqtDRdnYIDzrZfJnNBYDFKwJ7GfL
zD6eg9ioAWWPEwYV4nct4TgZF9cu2bRQeRU9JKS2AwO25jW/vls/fZRH2gn095shT4C5ILzpPd0Q
GpgrX6Ke+K5w5qltUjs0m38brb6rid00Q1RI604RLiiIeBJW1ApULp8dvO5uFWwJeRnbiLW53Eyx
9XAt9dfJahM8mr/FYDKki71nyoknsciplsRTXl/cyEp3E+5d0STMc9VEf43WyP0257LRwxgoIgm5
nrtDURDPwRxAE7m0kf4J9YRD1N+jAIHC1uvd7D9ofcAIOxxH9mBUTnkc38bG8yXrFjrwRiWgkz2X
t/o55EmBhPBAoX+9GcngDkCPImNjIIzmWNOM93rCK4ytRHa+cV8XGQsNvMXcmpFU61Ac0jdrCwX/
IofSVHBtS0Z9I0kPZsKraaflqIVjpg4FR/UKFovjcCvElhkcCG6TCHrtbkBmll5EpCbNP7B9VLU7
133A6XDQdV1/Y/ZJ91D7snh1DKbkcocUqRsAdlkWNmApD7wGDhbdFSOqxVgeTLhr0ZQB6iKThUmS
Jp+3/DqCk//p1r+RI10F0TzJXouHzddz2ci9jJNBb4KsmrRpSdzZI1xdzVs5hZc/vf47iCKKoK90
g7jkTrNSYRymFZgGPu407MU7jRRXJPVm/x9HPVIT2EHr65MqeeZRhbmxbOtuTV5Hxh5409eYtuWp
ZfzclYomhqYqKatr2OK3klogyDto+OgSdzfjqMNW6yQaGUTKQaJ49MmkEc2QNDtwhTTJDvFuccqE
wQ/MOPabxJ+9UaC7iTlhpNIp8mYJgtMo2zMFb7Daa/5ysIplqlr0QVSOgoZk0TYz452jq3T8TOvQ
kaL2HrVLpntdCySj+PFV5o9hPTH5aiqpwXpKeIWoa5LcfRLo1VntRSPt7NZE2MsAJ4qHsp0mDvqf
Q3KEPFkxDKut3CJ1XCGiFvIWj94HYTK3u4argbqSBvLiTIr/SJHrbeGxF19l+pPwHjUC+74QQucX
CLfDcIYn/SLi/1IyukagWyX/FRfwMzK4C+HyFSiTM8zwpE55/XvIr42DrdK57d0RNQ920siW6xao
yeVz+ND8wN8QrKfJWa6n/W5IcPogaqMehpeDyWc6TsgI5ftl+h3unZMN4+mUDxeD9q64t3Q9D6hd
sg6+oov13xMVZcHWUPNXRQ7PbnPR3f56vHHOOL8n32liqjve/ydq7xnoFkOzMgwifL+kn7fXZxgJ
T6G9hK1GOTjqnZz9tFKZt14j/Vjjqa/oo6vvijaRuKtMYyZ7LhouulH0NqoNqpMvv/lSeBDOCyC3
iG5sHi12cOOWMgFUk+O2dJE/Wl/DRQrkJMM/rAnVP8JYob7LIPoH13iRMs+Fp0xk7lSZ+GOfHvQZ
IkH1TVd4MFqeLKFMaNKVEHD+5xvqOjuzdpluV5uASVAvTn6uBB93lyqRyCedCtTYfZQLvJWgxHaj
73GRKyqczK+zv9z9oQwRYv6PHqwtXD9pI2aP1jBfn503W1WiaRv8/pnxCPStDBUwNuVQcp5BfI7V
bDxKcizZWIHGi2wftuOUJ9uJ6k620w5JDbkkgC/AVxN6EWRqMB7FbIGva17PK6GTf7Yjgn2UySbG
j2p17LNfyXnElg4OWhGtp1mC+UxtitYdArr19Cd9/JYWdCcUWecb6LQzqTVPRNXdfLOfnUyhE3QQ
aThwNn+hqNX+c0kXSF1Vy19NOq/nzY0mdoSQeHrW/9ghBnzGGc+vI/PbXwyHrT9QvZKpTxybj/qi
OazZJl+WcfV6mIWuz/CwVh5YV9AS65Gh9rkwiO9VO8kW6sm4wUtfCxShM1TYgCHfH7s66QHh+AA4
wxrRBNnCR50xYR/Q0f0LjZnNrmm/e78EZaPHXGlGf/Hyr5mOHZthhriRuE17Lz66kIS7zr4Cqq0A
kRmN341y/pAfJF46yCkRpWr/ps0xORDDGPjWcuL6OzomeN3M7kqEhAfKijiMr52B61f5M8MTZXBq
obk2/shNN/ZWGtnKR+jVMm+1LbK3U3dv70sKBtzFvWVIEWPZUeDvv9zVMJIdIXchKErK8E/bTxpo
lDLfnBt3+fbx0xLHWbF4fYiK8sps7KzN2lbGGAa7KVcdo/64KASkdXnPvVPyPCx1kvDLNWYiFfAf
FaipO9UlfkKyzyq22x4BUtb1oZP22mZ3ouRC/ksYvREQfLbnbyiNcU4uF8JzSZHoQXU8IAbpc6PM
YldNptizOIIhNyM9IvJjze/Yvkol0kmmMMsCbS2QEG1W0W9do3l/dkiRKNktT0ccBKwKMNENvs+U
2lcf0KY6oKIcWSO+vgzbgJg9YbaLk/FwQQw770QxeauS5lG0nmEYv8LrvVac0liGPgW7lM1A9k+e
C3oju1Vr4yB77NEh4Lwo38z0fYSxATWJN18SWl3uaKk0BDoEHz03NYVVvMgBtI4OVpyLpVrckUtK
fFY7Up8gczClEW8Do9c9FJTAeSZWdDRPDQwNP/1CQOIuFwG5lXlFCY02uxWzUHbrEHBJ7W+C7C3r
hWQO2t+xhK9UlEWZeNF/hfkCy6I6e+hti2FuWxxf3hoddThyFJJA7YcCxLiWJinDBu4Ne2dNlqpt
LvgpQt3FDEafp9P/ls8G4irFNFxEpYzkzy+a+XYBQZxn9e5Pygy+9Xj/qI/PNi1LOqaaifoPzgJZ
4L2gvorPDKbJ3W/Mc7PDhd7Fx8Mvz9DFQxXjKSdqHHqiASSOysBtAr3+oGYkCu7zt7LPtAfeu2/u
mHwCIC/KjYVMWMlgBJxBUi/tDsu2BlN+t734tYEqUv02qt6tBOs994eBt7mAsG5tyQbT9KXlySoB
FBHnWN7qWk+gqWfBp9U34L8+N93AUVXdCBwtHRcjkshwYkyo+ljHtPGDLPJ40cYeKvQTQVzBjC+E
1OJrklAy9Yc49NBwVmEU75FUHUdarjHUXmUaYd7usTeg+s6YvJpSRNxtkhgh2P5JfXYUUP3IEpe+
rrGP7gUvt8EpxzP9fAdtnQ44TRfZ2cxl45urSS7couQ+ntwqJ+4Ape+eGiy9u8yrHqUs5wnKNvSN
ozN1HYWCE+sSTTH9OwQ8CxjcPsrb/XoPWp7Eov7o9CNx14SBGVJtjmRskGYMby6HMtp2q9FJ2T/6
juyuK1zLSygtO+/uWLTWCs3MpfJIeJxoYW6fzgmev/U1UIuVpYQ4Aw8WpV/8gust1qd3k6+IaKJK
rHdxlXNFdkIjdax/xZthgg7Pqm5w6lRAPhfsPAwv3xiHUfB77JcdBRsZChJOkXJPaY28xZ8Th7tP
9262nVG7F31Kfb4+tO2qYRgwdx5hH9Mb3wgAJI5MLA1OI2TUDjIhBfPgOsntV6INXIyUrahhJfNT
p7GT8fHPbT+il5K/P1U3lI2/XfRbhm2xx/a9vGs1TTy/KEtdlk2jcnGfL7QP63DJAr8IxiyOcQ6k
cp41PxJrvSzw0R8fTPGo8oNyiZicjCB6xjrcrHEZoZUTgvGtUPylhtEfw+VMwQlB8Z76pOL6ERWU
Mr/awmEfgMb+ApeGm5wT9ahUHbDg1i2G/8vPXGK5CkXC8KtLEs/MAiEZIx7cUiMUcd27yD74Mtjy
AQNEQAJdLhhtCln3EUoR3rEkpUIwUwBgwjn/sznX2bxVTCTCGtnEZAwnApunVCJK9/DjZ4CKcwCV
BXuwkCfZ9MZu31bj/2o4AvoAtX2GadZRcCvt4e+6HLz8LPn8eeIqaLCEnrD8XHL1M7ujRRxwzq3J
L18EiE7HhVR99UtlZmkYQ2fRR1HIE5I+pQZVE0ww64WgzRbjrn7JKnI09wt6JIMuq8SYz/lFH4gp
0qNQqZ9pz8jXmarqOvRUsMmwb2FKQnj9vJxTop9MikUi0XAMFVLuicAdzVYztIQ2+Vj2ghb5zfsr
sDQ7ccv2HyAIMytVNYDF5S4f9mH7J+NmhEW1FVO+62QUtC90yCyzGXf/1l0R/JA5GmmjEIHqEB6B
9gcndNmlnPlXyss+KeFYK9CkmLcnrvIGH9/EBP0fu1K1U7tXks1zhDf3i+pGZxk34Zq8cYn+dAtZ
tM0p3DB9xSSmGeYnMnVmbN61/3jmr9j0KF4mrFVRLHhHP+N2/dCKuBdLZQnxQhE21+fiBeOsZr0+
a9ztZA3TT8GXoYCT7fWxpCvjmswZW0lcpLmlKnBxPsI8S9LnXwU0NkjtoPg22wiRML2UHmxbfYHy
x2PXPLpfkrHKIAx1F/ImY7+7nMd+KgrD9pWNJ9bctnLTagZIyyhiVE/vRJkyOaXrP5IqLjTbaEGd
evcJqOOpQxipmkTEH2Zfa+PWOFOq0AGT7SsILoYY8RMaQa65A36AlWyKzCM/2YSY/K5A5JIvwU/P
ifb2fkrKQLegFpJuhxzhSY+cKPKeVkixRxqZLC1tf0260VySPqL220chd3GkRPgORVGDXNEKcf06
hhnqt/GQhmK9Gi1usI+8Qi5eTP+GDzdFUGZtTyeh0uLyQwA2hHYHbRgy7yE7FHZrduc6HGlQCGpF
dBebMJQGrL6dPlxXJDrJCkJWTP6XjjEJo8toKs5LDY3UwXEeCdpB9CH2y7T+RQFCN9fkAqQkG3Ok
+kB2pXRxu+K2u4KmmNbO7wkc/gt5+Iw05By5I0uwIFYC8V78t/aDgSKKGU7wRDZmCLwOtjgHav3r
S3bn18/RCtzaD6JZc3KvvVxpnwCiBfBKOfesvU70EEI3+3PacF5snfncNggUl9XMVP6FmNv4PS7T
0i40XfRfFiix4fOXq84/gALJNvrkpC+m280c6yXkLRC07wS9FWBb3Y9R6SFoXIT/Ov80DgUzNsWV
YK1aThT0rQ1yIntKAnnyoyWRbUEio7wrvv62eCoRCY2EbJbGF8G53feTf5r2frESnye8hfLDWsId
W/e1Liv25Zc7b5OrtBSK2O0KhzR8gxapQnHYzhVzXsdMcac2jS8q4TAcSt3LGwmODZg1+3FaZF6V
DURkPagYvcuOw9i8VFo/WjFW0qGfGTG4TUnK/t5HKbTT0ouBlIK/rkkKwZnrfELGR7osTdLuwZwr
nIyzq7v8vMJY6gA9AF5FOxsm9Zg8Emdqzr5hko544CLHJ3gO6AMkKosjlAhllHxweFw2iEDpgdJW
s9anNGK49S1oBK2J1UiI+vX0mhmtCprI/kADGqxMStCoRBW3WyrWxx65C+r92hxwGCZ4DS5IFyba
FgulMQlQL3cOdNgZY2UXkkmGGTuXNBqsRHxJvpGF3KAH5CM8R8LLNz0iqNaJxuuCr0pq9KX/P4pW
M8xNST2aFQTlmAAu65z6QyAAY0m/7GKNQE7znctWmOtNokya3k61eFht6Zdhk0vuQWOnj9Xs86yO
6gQYilTo2K7HElBFE+FyPLiD8vANzdqiD4bnST+YC3Qa/kZebqihIQOVkHeHd6AUeDx/2GJE0q1E
aIUMlftXiWQduZTw7ntDRitopUB3ZN4iZ24GngJfRlCK1sL0GJFqDb7rHJydnt5z/j+5S6IXa1n/
i8Dl9Jy2TfB/NkV6BkNK/49BDyThyAFO9KSd+8pCKfN1EIElF2jk3M8CCWfvYgc1w2heKAMOzU0P
nsdcyNjB2YHQJRR48c0ZYpeobX2gew4TOkBXIxpZ3ElE3kvQ1SaQ2wWl0jAcirGtt0GTXKs4Rn+o
ZBQXKOF8qR/VY65fZJw8xATowdx+JHzhbsdwR7L+u8a4HmOQ6L2XKZO2RjoxcFiHpRDquj0Psbvk
4OgE7xel29u4zuF4fc2Sik8khWqqENftbID0DGmH/dk3kB4184QDYSKonCcNe95xDKjf7utoDSgo
DewMHo6rsoLHBN0PB9wxVG7go6wx/7cFPPJXZvTyIH3/D/3uZO6lHesLHDAT9KYZOSGwh685idWf
+nPzLcQ6jloEctlqo72tNpe9cgl8SGmiGJ8c7iqfOnhGM2gFGL+2p/4BUHV8RnD31ndff8XJrEvn
7AEsDUdHtncgI9eQB8LCbj8CHAcOrpnciNcwj+fnQcykarPlUG8rVnQRXEBJh4RiNvizCkZNxy1c
tBjrCqpo7l7ED/uPdvt9YDEKzqOZoaNRgODUy0ganFHnOYEwdAqRmCkrmVne+pPGfq9N4X3xXk08
UGyiv7ZRK9MZlVHWiJHyNws4j6BeDTsf6vomVtQzSEgDrBjHbysiqz6sgP+wdBm8FEi1cf1hq5AS
mgMhzrpLBg8EAlFWd1XzNpcXkJt5uVs3zEW3mPPXN21SwC5r3DC103VXZLet8wU/WqOwfA/tHWhh
6wXSguIqLgfAtP/ZP0pJ7/E5kZGWxhffqFNHj0zvfWXajz9NJ95Uaqar1Q9cCtm2KuDfSEzW3RVx
WIL3QcOGanbqVi2kS3sjRsSrWi6r6XpmdnID6PXXT6rOLhCVnPLsCZFzeoO0wlCtEWh25uyQLE29
3Svi2MXD7Pt3Yc1dVwiaF9/5pWddnThfkEoYK36pA/Flinhz+SncaCwZa/bKo1//oRBt640m2RIA
nPd1F3KHr62MKKxlxE3I/O2O7DMfBEG0iQQTah2WdFH4ELdA1p3stD5U+pTyC96+tYq4zEmUbDy7
Q5Gv4QLeKl+grSDYfUK59tbbJRxGA587ZPXPGQ3HAtVW0eRC5Xlk86Dv0d+kluCTJP5ONGhdaDFu
O17MmMOJN77jEwE0hX43I1+rqwB0/17EjmEkXuNkMGhPd1qv/ovRI0lTpD8Ax5D5evEgyDu3EMJz
/jgyueXhYxzwfq7skeToH+4pWcc5N4/sUGnUXgTrp5hJ/UpBy3hiZC54tt3eZS3RtxFEvR8aHCex
326EeE6tL4W89qCCs7PpgFYdhRyKJIWUAv6UZ7TcyrOhaID77OvqMZRIZ/881ASH2ValEvfQZTiz
a7ywK9006KSmXH7bD8tRTK1WCTtDYffer0QCYCT8ExbrXQzMKT9D1dfc1PS1sg5XXr6gYezmPKoK
fEpSiTtM/ekLYCfyn4JvZQfd+QQlcd2UPjCfs1m5TkWJ7ZVgWOcY7J8w71Oc9GF74AWPXNftAbMG
HsGNZcGEXk2gM70NGbsCyFJpqY8t62bnl82WWQPRpGClBH4fbRloMvMZnV3qZIsIkuVUXf/uD8U3
neqqWHyUUQT8A0vl6HM2ICz9KjNH/7ldrzIdFhJwDh1pXv5KgHelcwJqJEzxPgMMnrb2qIbd8eX5
3IEWU1U0aecJF5ycpCTL1Xig8E0lg/XH1Xc7YWY6nOxm9Pqlz1gr9PKc4rvwiuLsDwrtdlJymqe9
IcdvLDQUEamwEm9y1UD2uo1NxoMpd+c+/0uZ9z8ywDJ0FkPjFnMbBxrpt6L8gQDbsoQbTGnwTw13
SbCaWgtgIlkOvvmnyTWUXODB/IOwLnVu3PSrjIo9B9yiP873pQiSy1gHzp3XMvcc5fhuWBFLkB0W
YfOaWGq2iW8LNgZrIDSry/+QpbRwUeBTKJbtTQGaQPOYxFaxNB8qt2Upnl6uYPuJBQINpMLoFvJG
N5KyjMMlLk8tXJ1rm4cOZ7r/E6hJ5ZnOTcWdHYG4K6CpUyPJPPiFO9bDOYgnWXqaa1v/bLiB1hGg
4kYr3vZ6YgSyKVtRlJ1CvKVkSCZUyAYinYGw4D02Cd0xZ3W2E4fLxXfpp6sIUvP3zysgsa8ZJWkw
4heNZoGS30gJWCFOs4ilDhiUebyw1FhMIFPgGuy5euUsYAkw7u2eWal5H8CUjtL6c4638JXN5ifl
pN0keZhpZ+OhKV9fcdocRFliNii/VtvmimGUrurZxQJZUGZylJbYuYni1/um1ZxP569rJnLHOwnx
OJguMAqI2+5n+7PvF3P1XTBAd+d4kyoBVvGiO0xvdtgurT4BWiCs9Fpkem2cTDGz87TU2zHIc86M
UH7C9nCimt7APPxJveNsuWb4y37/SDaRW+kjYf4/RUlBHKKyiN3FuSavag4tLNx8fnamPgbtA3uZ
My3F95M0SZeQ9y87cuPK4X9viK2Bg7Fh5EoKSkdQBFuyJQk0T1GHXK6Za76xz92TBELuHkd0ef6b
abATZpSS2PYjCxRe4nBtbVWwMFH+EcChu/ORRqSwjdC3b+oVktHTe5nEtXoYSU5QVzETKEzQob4z
W+mIDOhNCDbiR4+IoZdlklZQAiO0OzztH2PbBFNq0KrscmhbENLIUqwRAtXvV6P82cN3Tu1aMoce
6oAiF//n56htrTVdFB6COOXbkKz0Y5IGE2dDxNBh1YRfLtUaYuPxDN+aKVL3aFbbvLGoqPbCjoiX
ZabtmbtymYwA/mo4hHbXSDnotzSQBc3qfujwljnWJPhyr4Je0mf6cugrA9143kKlKfuF7PMKz2VM
5VYKScjcxx2KZcZ0zw7jTeQv5UBQA+dmk6ufXJZXIKp2iTL+5ew1HRZGCgXmMD6lVu1WrHvC7Gke
7hQvyvw8DVmD+dolE2mkigRQ80uoNAaZs0MLDUyS/AYbgNlTCd4CBV2wPFTD/9at5JE7ADxSsz41
P6tJmIR942q9PdU2W0N5Qn5FSSNSh6jWgR1Zxyw8J7h4lfiM7N/S9PjXqgiYjdAp+CDtL1gW34M3
YKPkZIF7xVYpSkVdsF/U1fFGQ5WgT8VJITTb2cL0LWw5qstlevEJOvD8Rptn9k6DEf4NQYovgync
/zEqBTjGJ27TdLwntskdV87ObRZ5fC2exZyE0QpYiDpvIG1QXdw30MdNSA4BVcnRcRRr09JbZE28
VY5IUS9iwgxQbwdPP6c9XLiw2dC/dwaROGGHZBAMptJGbAjHds4GTe7zFl7HaaQWgm3+KC3K+GM/
izTIiUNzQwVVi20EqUqTJKmets9H4OM5lU8fG6uoHivo7tOL3FRWj9XHoxr2aX+Epnkt8hY9Tnr/
cNOwOmU0z1iQ8mgRZz5cuCxYdFrXQkOS96qK0faw2dDWtG3q+TtPhA3nYfOkUcSGMmnDpJTHKDJP
PfaazPULiVGZLyd2zSiMQGusQR8kwTeOx29BwA7S9AWuHOQcmA7haYQOwA4VUqJKKkIoY60D8Qlk
2R3g/niYnPvmy+UTSYd79TMFnTYks8bGZtLNzEG8EYtFeP615IqgyXkDxtc+R/CzEcFRJyUOWqV/
xuBi249ZEmrYewGTRfx/XMI9gdw2fqxxFgw89pL0r9jpEju4QxdhSsQBL1t3GOs7hPEZXBQF78VV
twimShNRUDA05MevJcEsbqoDA3FyymZes9z/xq+OJ+9xlpD0MjTpTPguWjOp+gASAhn2YfO5f3dC
iPaYVWcQyN5Y/nrfXzDUGflFwVdBrGbVdZJrJxpcT1CvT6Yc08CbL9xpfmc34YRMJclpS7FpUWy2
z9j6onPkihn3equtsJz3HFMNh/GhsLtYKp6cZZyx/EJpurS72NDNnoXr1R6jEqVTc23GkDNmcX2F
j6F4bPjhnQ2TkAXVV2wEX3E9I30mcT0zF2hP7Iw/DTCEspGoK5gz8cdf/CJbFo2L7xBFsrI9KTPV
CrbVIgsWnFTNyWkMUjCe+HB/UFEnh6CHHT/hOtAdXylRcMBlvPlU4vNwenUruKdmjht7qILFx73p
Qgc0eIs5bFVOD4giHQQ0nhXOA3fU0N9TSIGQvROF6hlRzfhem2ESWoUymAWQECVzL9m9Xqjtw4vZ
zyiS3Dk/BYX8fB573pYHegLOqmlXzhh51z9TtmZj9gDQPXSlGyd19LyU9rP8iqRf4s5q/wLQjae1
TY7/rJMnEdqjPpUVFT8TZdsYpBtoac78BHXLCNmHVyXONCw69fIY8+u8ksKcDLdF8JJZLRjOqIo1
hNA2a2Zf2yGb+U1ckqAADJw/Nta0vOZ4fCPJWL8oTefjQSLbN2Sfforw+unhAVJurLRN2wd637iF
dxGR5kpzwyR9w9qX7cX0AgUyJ0AV0vABm7ciKZondZvNrJJHJ2aflAZ3wsgtW51ru2CVLye8l613
vYERjzyBaZ26iJRWD+nUG93+4O6IyZdT9kZMpwVCFWgnhJEXJ1+LbYccdfB48lZNa6bAgGpgbbLQ
NET+Ba8Mm2LUeD1mHRGmHZEru/Y6ZwEGtft0yCO+hPvU9+yeA46PlL3z5I4K4QLOgqDnQzE76Tku
m+AwLiKxYh8AufTmpKLvwCAV1nLJyi4SJT6XeTtJ61EPruihgvBbk7wyUfcDMIroWgvTKY4jtZPc
sR8TEEs1XQgW5p2OSbRajo1UgS7UENwaNnf//SevWmcEBIOQgXqPi6N0Vra049OfYdJOEnT4tO5H
U1kHq4geiAwVAlSi9e0BlosigQrhJRaA243tLq2KPhFttU0w08qoYBQRA8eYTA1AeL/fPeL4sBF7
W2TOUD0TXoH0U78KVeM73EgERPAneYve2+APOTcdv2CcVLwgA5onV5y2wJqaUtsOrGePwDdyGcS1
SqRy5uobptyHSma2WA/rU1f4I5OOyMBXzjeSwC5hpIPaJ5hJrPA7p4PWOH9Fs8S6hjZELqzyswta
DGhDHhc6ADzCbL4lAFe+j6QLEky5omRr72q8HLGvG6y2U5viUDEGTrDVahJ6F1wLGDb0ESqkiOiG
eFA75s1rAK1P39m3WkY/ImtDX/K9/XPOv+PHaQ/twP8aPiwll4KfVQhKVP7GnDK3R2ZA0PQL2E18
2AWZx7Fgm3j8p24GzuDmxCgs6fIa2pCNOIziFpZBH8P+rGEhConw04ReGtc+L5yBXGf4OAUVfqnq
WhuanlPKSiVYAjzoulcxkF4rSQ/A+wr4k47x5akmHfd9q9Ce0LKZCH5VyxOOYKgqAEocZuzsIKO0
Essq+uiAG4rmZfwWKkEu/kDdf7t7coc4Zm0D1e0cnhQEVbTITLg4WurM5qmcInTvIDOXiHc8nlwZ
JJPpMr62oS63fU4/oXtK5B/+9+AAhpAqSvYZ1RagPHzWt/+5ZpcI4F3qQapkgLxdrDPteAnLF65A
yEe2FBPLVfth/p0GbPuEiUKTrBwZLwbJkWEfi5g7AzTtv544GG6Y2Fdrq5g7mlUGeNyttEvuCeRV
BgDr8wGrTXR6nrg//9WvB4F5fhHoD39pE9Wdp5N2tdba0FUMEASHx7sH+szRn81W6deGMr3dpw9d
/RHR18naHnEdHRhtbmNhn+SRhEhTmoV9GVHt5wV2lnedXVfJNtldetJ8opVTfHDJ8pk6QzKmVeVk
NxUJFFMkfVndAVVf20DdYIEo1IfGlb4cvrHnyMBVV7Uwq8Za0R6kEkZKoVpT+RgahgD27gb1UzCQ
8OVwE8cY2WnqYLdVG/SMDm2uzUDiu+5WSlTSQ9ggrlroQcfuVAStoQ8rzYhCLnKAYaT0hHJuckyK
LeIgz2VCRg8O0t9O7Kbv/Pgp72MbL5R/G9/ewdqmolgSJbF0/ipXl6qnpITZOuK9OvpBTC/pROXO
023b+34uRUQy/DBv0fQfOkcggPyEgZwnsMbM2mWkklXLtWFBaXQvhrToNrCn5iQvX40rDT8WjBjd
KaUnMz+3eyxNLpRl3gqm8CFEoD32km9pSHDzeyZYKYjJDikRoD6XbAQs40rncfzxPyj5wVJa/JCa
ok1iLGh5yoFRUq1LU3w+oMk7yMGQwocdu5GfSBWPwrIno2z6kVes7Lj3mpcZJy8WHGIfNU6F4FjJ
Elq8r+GBjbH1RF84wUXWGurJWyViv06TUcBYCckeIo36u8f5j6jl0mz4O/XzKLtQDDYb9K+6v/wa
oA3mqUj8ZPsvOjfAv/tbg0XnR3vapI0tVlpghBs/6GIUPgmCPnNqAO/n/FUiYEOvQhezDkh6NE+3
9NVn5tnj9SbhzLs+ly0TVVzo6QKyjS7J/6CqwTvq8VmoEIjbDXJOwnpNrvyirHWWiobrqSwXr4Cr
hu/C4eredO690cLRRiaSqKzjEJsHw97ssZ0imPtFdo14Ra7lV7i3YKu8dWPf+KRnSD0tOJWpuJrB
zdFhI4K3ay/wx9z2JgSOL2v3y5qFYlqRkvId2ZN9PbMJxwUpQKamJ2zB3a2Bw3O6STdycho8XqLf
LJJpk5Fsd3lJ0ihYZ03Hc49zeyCfYib0bDyxMDSMq0zRc7cUtYvjoLnHZbbOCjOKlWEf/7OM+Osw
Oc9yWCjzOHeAqnQVFc48XvGzhJjJXYAGJSUHnZp5XuVTZNUTIIIHd9tcoYrLWsnyKkqn3m4biZAo
fQhFn9JDdZc/nmWvA4UF6acQxLm7SvhQb83TmaVq4+CGDqUhIyxGypSEU7Xud6EIkADPD4pt+QAD
T+xzKcExh8adFzku+gejrt2i6UCVS0SGTiHCbHKzq4yjq7buKw4SHae0jDXhkFDWk5opMXbtIQKg
SQBSSDpTo9+nrxcMpWkzAcT5aN4m+D+hYno2msDuf8d1oenEIFW3JeHfG3e25KbQbsVUJqN7gKRx
DACfkKCY3YHX2Q/DwWl/+cYAfvgN1xyoxz3IZMVnhKmqdmQyTh4Fnsg7XZ6EX2VOBAOLLiz87XSS
Mii5cPsyYlb2K9yW3XiPXhv7g8xFvzlbvr9ehRNRa/Yp2uIe9vqgPocjK4t8+5QBbA5QXk/8YXm9
Mn76kCk3KY/MRWlhkQ6N7i7k7sCBX4YZtPp/KRraYfVJ3kuLwHhCFj1QSv5EPwK8vbbm08VuJcij
L91hXuQj0dPkop+NiV7YjG/RR93WzOWtMB76JfYDmGGmx1mk/jVe6KhRmqDtEI4tg7kVZau48qBY
XY7qie5YHmqqtTfE+v//QJiGr2S8YBLdsTmEl8i9ok6R2rkYiBaKQeHe/h173LmHOGs6K3zsiY11
e6c5AXw8QuXR/uARGZbtHWBi6jJoL5xMhMXc8hy80n22lguodVYC0g3BwoIx2JXCBzHhBlf5e7pI
YTf0CcNQvmfXphVrjc2lH0Zm5BLUx9gyrkY9Lpmgnndfls6LQI1m1jqCL3coCwSqCn5Jhldw16Gg
x8/LQkVxsXrRVhr1Jhfrm4oiMs19cdhLjFIxIEYE6+Q1K0eDajZerjgmJ/uaL1fSO+p/njtDB6P6
b8A4uf3Hyi2LWzmj6HYOreq+DeuA3Jpbu4tvr+4Ybdvfei9SZ0tk0fZuCj/Nx+5S1MNMAcwDFK+6
ASP1VPOhsFUHwDPZmUks9/eK+xagJngnRYsJcH+d5uk+kaBz5Wqn6/rC2H7xE+5EysIqC8LYqsR1
uHCLx0JD84Z1XJ4PvGO+a2YpfVNomhmn/Io81MiS5NwpUFlfr35dFRyDrI/qMuum9svIlsIB2aFy
5N0DIWo5x5eDdt/z83wx9RCDYPO7PKf6s/pOkdwEDWMoEBLBaGrP53OAbT8kxZdAor9ZTrpWEsp9
7moRKXOd1rSVdtqbwUpXiI5JFj/mleEpKmn6x9sX10ePQV0GPJ2/WuP9zJ95IVKTVapYzQb+OaYE
7NEnV4z9ofTTIpoIDGkKkBzzXANXH2vLzNLbCwdj6YqBsZn2TlNykoEqPXmzR995aYbryupZeW51
aWQmY8s7HuTl79ZU6FQfBtT7FeBO9AMNDBvMb4ahRhq682zGbeIpk7JrKXTRBnAyAcBJUdnBH6QA
fiY+hqr6K95jIM5BTh90y7VSuUXOFJVz0xdolJa7HSzrOW3eFlVYpouGdnHpKD761LTGx+B8dZeW
7GjRR/iJ2lOk5qDa03B48cQAabqi+6vm768KCihgsfssFNXZtUj+ip5+nes9XIrNMJ510gs5Ffi1
ra+W2w1fiH7dzjt17bz29zMVpdOtqoy0oLUBL4eG9Bjt9/27S4d3zfU6/3vSyN7L3BqKlKxT8PFM
LDUOdSNEbZpsthUDOMHq0fAqSIxb70NbuEaJEWzn9+VEWrHva+4vsJlRyOTiOGUmPc31G0MX0WE5
SWKwcFK7jUQVaDhsrYK2l9sm+JegYfrPxhjpnD+M9G9btYc6jICovZ/LtH+BvxGOgpQivF0ftkV4
ANwC6Ri3cE6FNVBS5Z+dolFrPMRHV14LESTz/j5Xs6jwU//4BOQoWVxu6wUREpJE2Kre6CCunfcw
3DfI4zdSVslD1CF9hgmwYIzMRsv7uUgYv5q7fnJgoHuWNALcTmLwXd2DS4df+Gh9Tgp6Ch0KgJEt
Vatf4em6XHk2Sl0zG7cP/hyIKnHScNhItiH9hhCga16SPiB07der4iEF3G6L0DAWxx4cJy6y6uP1
Z+jYO5GwB5udUgwBsOj82N3KS4Ixc18gtgqxNYEY0oBTWZuXpf906hJ1kDLgjeOYbN3gkLtt2hA8
3WiV5h3uRHO4lN+5546Erky4bCWm5r6+aIsxec5Z5LHk3AiIV/Z9sYvUpMLGzN2XbS0oID5d17qZ
xVJ8HqatnE9i++6i/b8eo2yJtDZk4yBvR9H32nsMzcLWXtk/soy+FHNxtGMiO6mK099HGRQLyjgb
9ym7+ZJ7mv50tSnLvzEwL0GfMQ0ISRxoIx6oKZYCN0ijxBF+ODo6HL1iWPw7I2tvHi7q5BfAiRyf
1D0dhI7ZX/xRMz+QhayskZ+jtgpn8NHgMx2ekPlidHpJcxcr+RcctzjDupGekGLsE7704teBa6MX
JH+D1VjYR0JPOdgYwSUVakRDvwJ07UJbvu9Gt+9al8agZV6dDdhdh+yc9AqH1RhHCInrPR/uI0Oi
9CwB+yJU2Z1Juhy9G77OWKA6whSF58Sg7uavmLAAiS+OJnZ/U4MIGehImL5is6ONCFD6O5N7wJBX
5umfMCoJRJt0jsWOWCJXYZHzAcPJWy369PfdpE7dmIVoH+PyuXTnZ7rXCtormrFU9PbmTlymgbqO
De1aJaUsVCaXVHVtntyhLgY2Cl7hImnho0zCBqCAiruJsO2+JPJAizQIhiGJE2Om/egI/Dj+8IhK
9wAo7PMtAy21yBwE058NyquiZQmZvU34b8F0XZrNpgaUAXmhWUpJYOncbuS/7Boy0tK8x9ElCtqf
qXi1OiQ7S9T13n50/um37/kdzvVf9sjB5UcICKmJLurbcuWWyb2L8i2o/RcaTDhTkvBnxaE9RsEg
/rWvWLKtVMP+bdKX319FRkh/RmtPkKsi5i9g+Dd7wBdZrw9jMqrPRgQmi8BvBXV2M1kx53gI6IWl
FtmbsOFvJlNKMAwEdeJtBzR02TEjqOqbpZZEGKcH5j0nXOGLvbfLKGcMf959+pKWXQUNmACLVvgY
MMSirm6juOvZTvRVnmGOe7hfugi+K/TqTtEo0PpfaYAA+irjTkfT4zF3ImjS4lFvTR1LY+ioHRFN
amGxJeSF53DTRnwdunqgsGV1JS2MnBEimOEmAM/uvteiiKopWjgHdDs2ENpEXC+5P2j63e7R1XQp
iqVVz0igGoIgylCVKiAe32SgQVgckc02fY5DtW/oq51RO8t9cNoFa/PZPY7YchjafmXs53wft6ff
SgEy2Se6KLBdeNmcWMbO/W9Donou+PdpUaASDaeXdgnQ5KHiaGxvXcB6K3w+rPN2Kw/Ql6HwX8tr
hW/ZL/a1kJcd505GqJ84hZULqRCb9LhfgzX/kBANDeQxNB7lcVD6m1jGSt/D9xJ8H5sJ7KL9sjh4
zRcnhOlHslIVKnM8aIjy8G75+ZmmGJ7jZhjNqX9UNoKivZ0mgKs7eLcDlOFlyBv8wJDus2cmfbjB
P0DjD0tqUWznuM/GBh0r7OPE0cdseZq9+8593lVqknV6C2iJb9Z/OCEEwW/PZsoAx5c5XlOou8Td
JPjkS4ndcACiq80OMTjoaFXTWsCFVHHgbfRFBG06P5AyUldQUw5Jk5eoTD7SzyPk/OiCBoNrZ6fH
c+joPcvhtjR67irNImGFw8OatdRe3RY90tkS8Gara1MgYymEcUiVX5sKKExf7quXwG/qLoYpJPng
aBx3mZoR3IO5s5wcTyVlARTRMZhSyxUNAb17Pk/Mrf2mqOW1g69hO5JjMhi6yTvzgLOw8ABLhTLI
38V5SGH+Yu+LfZSenWQqv9AUYbVo60dJPGNrF0IblwR7Kzxz8fi8azwNyq4BNRNLChsAQoc7aZ03
SKLMhpO6+7x7nrfkbIKSKYmRUKyWKHXR+XASfWJIPWp3Eape2s5133rLD8YWwdVCMAFKXStTSq3l
e7Sxs33p4m10GCalK05o2/uTuqd73aYEiTsoYkZkoLCgBLV3ySyml1C1mqWkSdjj15kTeyNC0KH8
bdQ8Vsx2y8RKqcXlHutpPsVzinVVDDVdSVup2ZGsdL5JZAXIQW7LCUCt3az0UD7Hw8w2C+D8AE2F
sfqna3RGXU6W4jCiQ4+q9Uhoq21AfKdNo+d1Ry5zFso6xQAoNigWJABiPKFpFvpoxGhEIW0AHx9O
pGeXukbRr1ik1gAtEbzemmbLb9wsXBYkg6atoPt9NtVHMGRCLGdk4PyK+XHMCEcfMqZbkjkP3v8+
or5mJdaDWZAaY2G8oIgZ8HJdoZQPsd3yXQD406DNal1tnnvI5x8/zVEG/AJi1J1CShwBA1251q3k
/KnhlS2Nf4ymydpYIN99Rgibj2JToCUaQv8WO6DScMpAnKWoQTqgJWVDt2T1JPF5joV8JP3e3lju
AltyyYs2zzrZSJ0NH4n2jF0nqZGjvGjUPkC5gXio9AfZ3BiOMm9xiLsQDCqfO6qGg0tOiFDUluUD
jgzuk2djMRlJqoeiV+oG9mN456g1Hm0W1/TfG/LH0P53ZxL+ErnZH5Xid5mVND7KaVNJni87daVq
+3Z/8/FCvXSi1F86mmLWBmf+kDGLUZgcExNnYGRTbSde1Xlj/GXONcvGJ5dvaWded8WnO6WNQY2m
J7iHiH891UuIKf9PPblTKmlaGub0sPw8MoZo1BTWJz2TdhWIps51wR9foUqTXLolpu9KlmrpLqqW
lvHkrlLbxQXO+f4Y5VHqMBTsDE/G4TkL4MRMR+vPFkJtYsa8alt9tXGEMBpr5e3p5Ne57nfYiltd
a/eQusk+8dcPBVSJmMwCdaeddMo7qZBlwLHDP5TeRsUGtUYkgcZClnwoUxrDPGvlsJr5sTc/tGKO
yO1DVBiKJurAlvsDyBCCKvc12aMfFDyMBlseWNbaHRb3ZxHMN48+ZQmtxo0pHRvbw8x9PkZd/9IL
fMQuZsq1Q6pBrGJeKp+VvMnPu4Y1jjkpP8BjK/RsRSLBOrN4cWpc3HXxSea8827MnsLo/+l9vhqM
MJPUus+riDDitVDwGYIw0DvTFVHXwVxbyY9Q7uN26LI+u/T7dIK8cBTPN43taB3WWDF9pEVyP3Dh
0lFTaY5R1g7ylX4dOLFnZTOR6cYROVs5RuxVZPwp7qAGvD6KRdNyXtAi0DmOZIm9imH3RkV5W+gi
APTOJ0F0G/IvZoPa5TjodzvlUz+B+bxzbx3nUv/ZqUDLfsZ/14ck5UTASK4HOzq8oHqn2elb+H/6
YmcTQNaHnrhuVXsH95+6sciW74dx21/M5jcV0/GcdiKAd+BC2z2PP55KgAz8Woua7Xw9RY9nd3D5
qzUwtlgdLk+e+U1cOWH8SAfiVaGCCr7Qy1VICa5AoIdsfh5pzbmejfbjyXXZzEXNxUxzo/4YHlbA
wzFjo8jK+o+6LpUB0Exg8THocbvg520lxEM3YNqlqZMul2l8jRfRRYk2GbhKKZmjTNpSIx+FJHG7
S3PM8WWHQQR7K7dtSqJM8nvujgqJrcuRY/tPQUtrQzoDKjRXrArrzv/SkXVsUJOd1VJFf9jxyKEC
F84026WU0/lOUGRw3jIbo4BEMSBt3FXax5G7ANlld2AK9U0/ya+J9AeXPFZ0VmaX/pwu5UKWRf3u
8ukX/9zCDziNIf/Sn2eldnbORDqVr/j+UTcx+yVUbb/I5BnBoBvhs/8Bp1j9HaOXoXkEDI3GwL2p
YPWkQV0W3s4BXylN6gcP0l+Lo1f6QQr1UKbix9qTgTxxlw/cXfnmmWhqTzjwF7erKCcw5PCadR1R
lQt1mFbLzgXHwyoMmtv+ClD1WExf/BpC9/gzS/2H9mhYzntFADYLN4OsL1qQeo9fv8iPTLh4VGDe
iiFjqt3lDqrqYdCVzx0vw8nKh0LybPuuZw/4Bba84Urv5Y/J51woXp1xpBa5DaAySFZTc+vjtG+8
mmSwMIC2afpjpVekaLx8254jowHH3dPGAL8QIuyL5W9DXCs=
`protect end_protected
