`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gVAb7iugiIRokdgiAVsXuQttYQHqh6d2Rg6GZfYvBIYni5qyzGMo5rUKYL/V8o53juKbg3Ak9MUG
+Zv5ERJJew==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EP6weDZrxIgPhe6B0gdYrbV0D4/lrcwILBLdzTECu+V/VdbEeHfTm3gfAXAgMLwuOzpKZQ2hitOi
e8En7V/kVql9zVI70+Rl/Xxx1+My32c9zLFDaidmibjytxCXMPQHIowOrsuz6u+GzJo1idJqk2wD
NgPfzijCZJTZAPh7reQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
yiJxoJqn9O4FkkN33BSBKDY4Z8AECfTIe7+v7QBitxOiT5eP13VU5kP2mMn4+tJhfOMdrmJTtrda
3OWjYw1v0AiQWiF8CXYetkeBPIzDP76xpnCCYEJbdgh9RjXACEWpR7+HFSIDZb1sTmhS9psfSmGj
579jIpjzI8MVhlLUoU1gvSDMXWsQsEsOYZWZMQkgxAZVA+b1ZVbdA//tUYE4upskQbvxWSAsxhHo
i/lC5igkclkV8S2/zzDuWCmLOiR2WE46P40mw+OYxCRDEbnFNLtKBiCAQUgYy0jaTM6fFzlxjx7n
rLA55iEXDhBLbZBMJlmcO0xqMYw20ueNm1q0OA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HUlZ/vjCyNj6Lg6SqAHrP6sS3/aoFAvuiAa5co7cL1O50M7zerCzvsXnPgrEFNRBJWlcATW+aM28
f2fZbsslFAseXDe8iAPMpeOPJxgHbe5mBk/JnALUBS4HF/WbPpkU+bRrZJ+Qlr7HzSsxXiGLLmMG
5vYmMZ8VVDmNoc6baDR7rt1N7vunO3RMUYKj5xr7+5iXP3tjXrnre+ja2gc3lYu9lIvoI8FTbDkA
gdmSD0bPlJwyvw/E2o4/xxTaoeVqso8+lnrZtksqItQA3QWPqu9fypgc/3zrZLWAx8KVk9H9quxe
uMLSE2ppmckotn02wMBQiRQWTE+zf0SHz0qZTw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IhbhSOC/mglN7nLRBAuGON8aX15xpKkqAhqjzcWZdjIVEV7Gw3F9IYWlTKiwNkV1BmYlwEYmaxjT
PI+s96VkmsdXCYV6DJcfJFFNxWOBplnQX16RUm05474sxYsYSrwbLXGRtGCQe/jOYGz1urfBcPEz
0RZC1XlbuwihHvuyWsY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S8r0uPAGnwkhC2v5KBlF07j3Un+1pXM0dreIQCvqRXwzIuirp9Fg6eHD8I5a6CD9Xrl4geYvYPjh
duyNW8G+Ae8+PMqck9tXSgZGwcnBTyoWzkeVMfLWIJ+ONkQCHy2bMCDHIAqsk2tRjCakRCOhQqOx
Eh14JZXr3wPdAnB3X4s18HRc7jsnM1jQITyO8pOsElusxfdRpQiAotN7B4ptyG7qA0cAzo02/OyU
48y4WTKg5dZBal9UoV1MYyl6qO00bFocF4shFCIs9exsAKiAKC7cO8n/W9ifbPd0GT8XrokRLA4r
bIjWRHa0ladRVspTRoGYmieDqMH/b9Q6P0X0IA==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ksrg1yMamjhmeTg+uCiyJ3+Kfd4xyYwxLo5/CmGm4mRkJZDMjdBNJ7Og7Yp1HqGdh98HfsQohDll
ZXP+L3Vq3bEx1LMDpeZl5fsYSQKsvomnSzPnN/w0aBcGMzj4sD9yl1tyCp6rH3GFwUWMnZhiB34A
KEkt58iCpV67V7X3p0nXW0NPXkTzuN/pR08bNzXN8h8xRSPX6gmVvuGjlD3ydyTMv7HCmTmz3zgn
KiJtMBoaF2wyj/JtjtOoAPMblMF3w+gNJh3vZnnnHOEw21JQmPNMOGQA0izgWHijz1NUFcic4jFC
Wnjp6UoD2M/+JZLTrMuF8YCGKCEQeB/BVoUTKA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
v1MP4YPumZf9lMShN8qm1ipU4eyKoQMQ4Tn+Bo9ZV0+HuOqWo8QpDSu6Iq0tXJTj3IUCqvcHx76B
ULMmeWZjXaSitXt6nGcs5kxU4wse+TwCRyaDXNhpOQRTTCxCCLUPKUJH7N1eu3bknqL1g/qJzhbS
FDnTT+48GEMqbdFST1TE9DkOMTc/NGSLHYY9Zvf4xW8q40+jE6kKLpqd5DrvPzyVxoSDtwjbpSmY
6tqB7MulmbrnokyNJIQrqiyNy6+jm76tJyyQoiLK3lsH6tz7YrQo86RljUkGrV3lNldXzmZx44xc
BbnCFd/sPOtRoGkNCSRj9hLCJeRyUSmE8wRiTA==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ad+97BYKefNZtaX2KFNRZSF5Pydk3vr4xnGBXMo8/dX1cCjcqEWT4cAZ6JgL9ZjkvFnCDfMgk/gv
K45zBGl/3qjkmDN2roqY86P/MiGWfYZssOhqskepkw6t8q68rCJZzTvJ1a7ucpHF1t+hUONerOgs
XTfDNk8bYnliWa8724P92F21XWMSXFYfCnu1L5aX7a9HvIZhmgpjnxv78QYB7RKKGWilyIFxFWA9
gkmKzhPINdL94gfVVuSKT5VxX3H2GCIRTe9AC/DnebDUiVWA5f3oyH2ieL1noPzZkQZAxh870nNH
sDAtytYueWqIbrApjiTC2Z3VIkS9PoA0xSezkg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 566368)
`protect data_block
rOme5njgtdIzPRBUhRaFLnUkZpIGm31DZvLC4ghCtYmA3ScUhZD/euqvtwhy8v6TT/dNbUe2SrPR
+g3Btb5O8j7FL00yermVu3mNdxVsrRfCHrehs0FZClbYAYD4okLdwWiq8FXVq2fDOWkGAxuDT0Na
OeuIKdqbOBamEbx/VDb1MzFiKT0yIYwNJSDbeAPQfVyHRzQL4d2KyBjlA9YE7ShdvyVeINaQ0wem
ZNEXTCDwu4PT64wNn2cianS9ZzK2+Ju7XgAjyWyZ7tBfZnnP0jv03uokC2Qnquyuh1IzWcZRpyVA
pRHwERbNMuKTmbytEfrRf3lfV5uDNP92jRoayoGECA8wsPGuGCGVrvsa1OobQXyetyZ/NqUB2l8J
0pop/OPAMSHvSfV6UcZFmylw6zIKRKGEXUsbsy01+1fv+2HGM6yfBBFTYnis2chBSiKGyR8uWv+W
AI5V6NVq97oPbNj7whaDqTaXdWGz4+/GwDktCfoS451hRSQPQQWAR5LwA6f1kDPMk+yrYf17dHOQ
dI69iSeTh1U0Gi69OWpUJq1z4/WD8LvMsrlcecIl5p8M5elUoTLMGep0f0U7vGB9VHSynBTU+k/F
nN9NSzP3wzBQiFlPtHfjpkNTtb0YNormnHr/r7QEfxrQoCCpsqS/fFnMT47lbYEJZyAKRjJE1AsB
kgcQ42TBoATP+Uco+kH3JV5e1LS+BaYof6icp3apky2XSWGQTx69zp284npRaomk9nkd/u/DfbJJ
D4N9jpSC2kFcws7tMrymEbN2grnR3VofaXsMibYOUyS6lvldioZy6zZBCI3gpls1fXhqmOKCUthY
liAMSQiw9cPlA/RF9zLjjdW7s8YOjifWS8Cbota47watwC2jtTfJG8/0VyjRQY9/FHykMkcVAWYe
lcKmO823OaXlTb7apjksE06JPChOUW3JVCFmXCFPmXiwgyDj01UTdhxFKGt12T8Cza1Rfpmr+GGe
1cxwh4eaHZ9DnZM/Oqa6bCsCprxdn2Y9ScmCdePgwYWEldgM00f8VoYBbj0Kgr1erz50O/zlZPKr
HRSRulJdReKGKxBG0un6Mv3dbbsi6KvF+wRPBdP31wNxJBHvIJClN6OpQ4n1YmE8mn24C5sKceBJ
4kuxGtdVL4kQaAp/a3afXFpjYMfXp38/txj74FXqnf1Vb4dG7V6liP4SztMAvGoSWGkvo1zazdo6
HKnqc/scfD7mb7+j4Wz+aE31XCGwKUuPlcHL3oU4/+V9TboYrHZad9ro8leigZycYWoykYulH1Pe
noxN+Lz4GE7S6vhf5DwM/ZRFNq1y6FioiXBh1YtXsIy7wy1w09XLq/nEPd6RIWqDnak3YJ98p8/R
9ctLHZhyyCRV7YnyZTU2uhyGn7efvWNM0B7c9can3LdLBteW6oHDvp7r4x8cIhcABaMjQjK5QydK
83oqeSoalLF00WT99RvZaCz6oxbYzqmIgPSUjNS9jJUybC5i9njJitHvPiiNd2N7nkr3CoNtfF59
qFbd/0LuTE4Zmf/EPcbvDLSYnobKzbdvBfgzZcfpIHyLTvpSLuD+F1Dye353ULCBQ2p/XIjmBcXZ
+mZUJlK8EG1GmpKwFgnu/BpZC3P4iAHxrRLpbTrVBcd24US6okia6jMyAJsJATjmM+8/YbmJvUxU
zkXFDmkVcXdMQvx0Lci4PuFBRa8X09b39xMSZ8ZadOKdYVs27Elqj8zC35KTymcnpiS1YS/lFM9q
S/UX3BVXcyHT2PUSMQI/XgMxq5NCoYm1XQPjYs7fr0Cal0NPg3dTDvrZJ9fUEOKTKVY22YefZQPD
Ej01Al34qqnRiSWXvJIwoFZ8Qu+xEEu3kergpqr+I+s8NHpADnFR+hobzEYIfmoQhe7XCIipqljU
V2FU7eKCEGE+1E00xJFnYzjs0ufrG32ojv87ZBCKZC8LHmub2gTJfEV3v3QT7rJWSuIjnOpVbI3f
d9wQkFW97NNaCBnYaiCPjlHHJgPn3bTN8mlY1lIZrijR2bMpars6ZWhpEt+s8t56a6kMkHtNsh0B
Y8+Hq/pgpJ5nJF1dNx59Q3D4Op66l37ULB3BveGUVaT9vE1PoHZZe2bmdnjkViw/t0kO97YIPd00
la9iPaOHXqMiPCCPIISXBENy9om5W6P0QjtsLF7eSHJ/rOoJWd9Eyp0huNHg0iIzc1Dd4Ak90DMf
/x+tIiSU+LGL1bM3bGQajvy9SmVhipSJCUYu9HSInuPey0MmTB0r4bUM1C4iDMGoxQwMNiXndsll
ziZUuuM0rsEliRmoN/qynrUJ1sGgr0Wxre3M6E+aeZUJyfA2fEXv98gr/n4U5i+gCfTG2KLVofzQ
swiSVdP2FN31FjgOS0vIIPYE998g4qmmhRbw0lWYRsD3A2nsuYKN/y2aGPCD9wK5kcNUqf8I40NV
eOVWb526qvE6Z9pAAkAmBcdKWWFmMwMETXZ1tJ6heJGuQyfmCiYotJrTDV+jTiBIOdQW4eDn9yPA
z6FuvYn5xhvIO7Axv7KN9m+duycmsbuCZvBgJn76lnJ0e03nOxl0cfZY/OXzcD5U1sBTvzrh5X6Z
X03yqcuO4CtjiCGgIOryXiWUN5khkZscso84qgIYIDo0Lg54vTbeObbtu6+QAw1xL0o7q7+bzvJA
Iyx9UHHjw8+IhzhnoKPym4m07WXxcqSXcLUdpo1hLQDkONotenvB58rfzj7u6y1weA8s1fb8HLi4
15A+2rU/cRz3CdlBqVPUIJtRZie2pTd8NhEm8WuNoFInMdGNlAeXebskrQB5bD2aqW7SdcbOXkZk
CAuFveRaDZwWh3b/Ijt/UDpDZ02Ieu73ZDMwypNXIxSyEgoSgrksZ3rMSnl4VN1jcrjb+7/SHmCT
CdfVQRbGw3pTwnibZYuVpHsVp0epOiKc3ZXZC3qSD2t94ba/iIyT5rut9JMdV0nXkEdIRi6haBUl
Fgg7lquyfy0YYMbwkvTjO9pd63V0/C4welfeCZ2xF+ocQdcxmMzZ8P5wWnD4QEw7T+bQ0dKtY+KM
AsnkuI5IHDxYP9vFhGlIgVSadjkMgeq5NaUoGcQDwnmLJkQoB8Y0G7v0VIcyyNCKIr4Sh1o1n6Cv
bP2uo8n8cccWDH6ovln29LR+PSLKxnaVIc/9UIN8gtcgtr5WXuoKO20AK+91flNCBlJMjES4XZ5K
mgfbyiW0e/YYQtmRiNAiqU5gGMIT9eesVZfNkO1c1iRI7HG6txmy3txSmAhAPpHkI7GHpmvn8kT2
7x/nH0wvV6si/7t9xbg6g5Fwu1YLWxCYPqdiEtm2stjD2PA5OqSi5uTouYJp82io0c+E1PmBVkHU
hrSiV88ZMczBkBovIhTZmqz4F3DOOjvwoNWh0qsoGRamg1vQzMZk9M8BcubtWSQ5fe4d22TojBu6
yQHpY2+QMgitVp7bR87dTCo7jJz2HWV9vT81MLQa0vl8hvHQvYnx6qKAW+Uqc94LOrDsOsOIufY4
VI+vBOidarEbX82BKCRJm870i5i8tuUQYdkiTM/YKrALgM6/l8PrY2LSctmVFb7eF/gGmLK3Ivqw
jULBm7T7vjs2v0RBe5YlWCD/0d8MZX9QliaxexZcbpWi2nmYHWczj+N1x67A9L6+9TwqlMsq0SJ8
qe4hzqxJSKGOC+1SvUwtBcsNzRpYCICZJ32l9p4idYfx7QI0FwDflELjC8hgvALt/bxgxontdpxc
OmUFfOZjpdVL68NzmkuCHMOBmd6FQ6lvlkYKxGC9NBQVPfePJnfXFoFlQoC93AA+n+rcjN1Ct5t1
8tkZ14U8phNqYy4LHWwl0b7+BNOk4ngjFjvqXeBNrparTOGMHwmnTo4krmCxq8QvwguESg4HFGbs
wIEGcQ0wx8Ffg9z4zGseFn2I0NzqvRgwUoFpDSV/sk+/r4y4R38fpSJfxmFoF9l0VmCHH2e7OTTd
X3HH82zQmfEpu9Ib1cnL0+g6h6ZRl0wikvl0jNeOMDRt2Cw4wQuRSDgW72iMT6q3O8CyMFhmKM2Q
+0lAtxWUiKU3DWBFVHPhfnt3ibuUX0o0j/kC8yeCHryqfekBZL5QNilhPLYmLqhftMIbNvw+Hcyz
r0Y0FmMZzm4OfzssqoMiJvW2FCAHZGRzRL/VB/yjTAyzGHoTmAC3ZRm95jRoyTY1u90VACf/ZcvJ
eLwmQxITGlOPm5tyL8tQrTBHgYaioxlVlp2cqWlnPSFpZ2wJD/WO4/0ERyg0XAS7NnoIYFybgfZ1
VlDsgkVnvdBuh/wI4ZP+iYMQBCWuzwhEvimnAAg1ByubP50kuMbfNXRxtZsETUYsyeTtOBPz9q+0
iYhzm15vygaqCoouwwVrKcAIo9ZSi7N8mHEMadoaBdnIchLANo2pA/aSfEgvoBkak6r11ySoQM+p
RlVUBwBpq+T//1L9OjJzGCmtv2clkwOxV7z7+cOglCHG9jgPQpO9csfSQAnzVUCkZI8mEupRJrWb
KdC7uOKDQEzoLWegFy5mFU6gN3YqzgNoiiWHA2mV4tPtCZdI+JGfblVbrXVsg4xSCTH38RW6AnNO
xNzSNugJ0i2d/z1ryWZ+egqt4NIJ4JDGXZRJNtVXKph19R15NbZl37yQtVQeYh6xl96+DF/udCQg
YG1EGAChf+Pi4rMBNWHZHhnSPP68MgZ9/g3rMYHU6w2qiOZJUZsbmzVHbEEfsFoRo+hvlWFgJlCs
AAw2MJ1gxg1STUEkH1j0p7lPU3yWJ9QY/D3/Xx6ZPjbv2QRUYFpRw60ibfA7HWaHCjyqS3QQ4IV+
ngtYZbonR1mRAyk9k0pJIajS3dHNQ5p8uAdFHj5js8bKzNXQ7/K1ERbMT6JtSuiM6ju3zPC+KUi3
CxpYOmC9+6yG8Mc4gkAu0lCebT/3l7PS1XITPn4kkmF4BtfHdxWzo8CbGw2J9hMKPv63TPyKqa9j
7Umx48n2VfqMpSN05hs/+jRwlpnPiOeAaqn82YS4gcJTJrCopuSaAZUlyipQ1OUre1cy7Un0IUNN
E2CJwZEMj8IpjcyT0Ya2NASj6Aup2aR6QWWbPACdFfA8Pr9pKcAnk4BHLcDyYuU2m0kOtVpCg5z4
gOAdmusV3svWKT/LF/IczDWQmYpsbDqN2IJgQieSwzKOachGYnAdL0g3pZi72I2qximDAa2MqyEK
13rtzRFzJuWgOJ1/z1wEEXCwsQaegar/AR/Eme4KmkcNGP5D4CRb/Wvj1IvMmGkqsBlm7jK6By5U
QhBjjCU7TuTujt6ZmlNILNmrCBswjkxFrhyAIBqMxv5k+6/N4S8X35R9buG2kpeWxzZemzQQ4pXv
uGtTExyA8gSeubU7/Jb2WmlUo7g9ahXqV0ZTxqjVK88n+m+MN6QaYhrO7oICQY0OPl/NPmN8hYt7
+hybAyIZdNLhGXMnFwtiaNVEYfrdhi52MmSy51IBTJpw1m84CF6R+bUMZYPbQ9rw812wKLdroyDn
wY9i9sJVDTn11ySUHowcRLspvGcKXV7qSZ8sBRExh1dfd7xg7nzw8MB0aMXXWiS1OfFTJIJyBEaR
iM8d88PQNwpv3DLREwBIKua5t6NhodQQswVoy7ELzsJKV1sKoa3G8O1KrKfUFOjcr8ssoMEcTEf9
v+LOp+QHr+J+h7rJJKBfHh7Jx0spt0USseB4nLBJ18ST51CZAyRNiIu5OXKuQh8Y4adwA1UGCAtz
XLts+xBA5zCwVuIa8lNKM7BHAHyiwR4gxevSijqI8QLzFuosAa5pL+mvHxXPzszgkT7C+D1eQhcG
2suF1eUM4GNnVTsE7/zrFTmgLw8GR3U3274gZJTVOVcyDjwfTboBGlT7ODpFLOqloRyIqcGxjQs4
U4Ms/Hgz/gllI1QIh3HzvO39yFN4wDjBjK1N/sPX8PxE/vOJAtmvJhdOo1/wA/agQQ/paeCSyAhg
fT/AIs0xba8fX+4rDYIaq+IyMhL+CDMXMWGQq7VbYYjIHShdTb8GWzfQx7xRKpahtFabMVi0m4Fs
AsHpUG38uLRLeSzpo9SmDnms9lQ9y/5G3HWG5wUA0hGqeO19AXm+c3X3sln6Jt+GtXS3kzikL/5w
oo4G3QLmQGrKplYhSIH0DfCcoCt47BXULe5uYwH42/HzoOvvdiX62ZXGyHyqqyuTZtIxFkA17vkP
xi2lysAuXC4GiXc8OpRfOa4p/mkCOclzEeNKsNooeuvbhVot6EqD8uwLLpyePyjfcHoXcG7vgOBc
uQdaLf88xU7SCmWAwz6z/mpeXul3ZHzk+XcmomE1cdYD85xzcY4t8znnKxSXSttWqIMBNRAofOOc
0aTXQzC0NXOL8OdfZz6fSlSKcAmq3m7T19N1K16fdp8zAPWgWyHkZkUeN+fKTQbZlTi3ritxYuKY
Ab5PC2fIpsTe16sISYYZkH48EPGZkJh87mlkZKKC707tvPyLQRCRTNf8gFY57N4dknJzRF58IcRk
qbWimaQkoX6SX1ft3fX5GL+Kh3NTwVvhRSHkQCM+8Xf3p1Kqa3D4p9Is89xEPgjjExhvr9NQxk7g
lyyQCDEl0RLNnJf63inu9XYqiHrdFKx07w9pkSvguGempOvddSEZHeQ7s1K20e+bOWnIktMU4QWa
WcefLqig/W2Y8BZNcaZ+/eHRpTl6W/R/vpm3PCynns8eX4Vg0hxbGpLyLY8zVmSzb+9Mh8fNv4Gt
XkXYz+oWAlGKNCrsgl2K8fDwYGk7srlf5/70ClLg2hzmc1cDA6djwalB7c828FeP9GHlFnSCX8uC
/Yq+zBLlfb0XbPrbRVqNKR8Z3i7ph8LQl8AISsVbtX7aifw1UPz15NSgrdx6iOjUKoRrK8pvRxmM
Q3IVywkpO7P1CWyL1UCzS2qS3QB6Tc/PyXGo6XVhwNphKbNv1TYejlxHWRMuIDsUvrFdFEBy88u2
tgMbS3snY5RmYOn8Z/dUG0bB8BZC6WhJNcygmN7WSSRhSOTQtyILfgFW/MC+rx/SoK4uqAhrGGiV
AxuzmSlHHh4FR9vcDhfxi1kkAV2VFi24Q2/6jj9pXRmKdPtgYvvS7IIedfZAR9+p8WHxPuDvSHn5
xZxrIxGHivY13Tv+eQzoOoKd5DM4rP2zLmKqNUuKA+I94lSM4sZmEhszi3K4K/5OxSzwOp/dExTV
zmyQrSEEjUVWHRU8YpuGjLccsY/Ks0VmKjGE4Nw+2pSfgFc86eMqGWbIK33xb/PrsIdVL7Hv3kSr
hcWqYElhMWpMTQCIbFjEqFW0F5jwPFV75Ho234d5m3V17iq5e/YppgybcgqrygDMDLSK6rafBCJq
iPj+b8Iy1QkOlbSmz9glHG9llQHFPnkmm5HXlGRO0iqvBlnSPI1Inb+/K8pk/+56Muao6+9331ku
jV0Hr/Q8OVduKK8aG2klVqEtqN/R/IWRHyD4M9bUF/SlXOj/aZC3ec0dwlR41AT6O1wuG11jNxza
PXxWEvxsiXg8vQpm50GNT9GcNTpVQTt8ShBwEAWBfCKZRk4d8azPDB7sSV64Hw3Rjv7QSE0NUUG6
1mt/0JxmXZtMZV5EsUNJj9sWCZVyz+wIpjdfc/5WqXFs5pGOfh7ZmVOBmbKQJVSmQyDaAfhhKsgG
smmVOrJUmDKo4l9tffNJsVGcg9L5Muz09D3tU3JJX6NIjatSGo/3sIDt96+U1tksj7p8j7XKRcu0
1rqrP6GfWcpTS7pUUQZApoK+EI9ICpAeGPDrdaEJR906XtjUJ9qCpn/ByjVuWPLxFOcOqG6zFo7K
fsHA92SIe7ip/TyLHvhoRvxr/LZ1HIBlGE2iOHAtXdCO9kSNEBYgIdBKd276OwZYobgcyueDZ8VE
nh41TJIoNcV4R8A4qpBmoMoudxx1Si/h6j9mC7kuzYzLiuar73m45L4GwO8uU44d52hdfX91M7eS
ezB2Bb3vllubNgaSTYO7Dj3OMl6sZU5OQJTCaShuHRLqGYTacggFFjrQJg8VQ2mBhz4SPZbYTzj0
PhecA5xTXnWYl60weKwH48DjqeMOgQGGOEgzLAjWFsiiRDVQChZTiK0VXhmi8/RZHmwsQBzZtU8l
u68vEjKWswfPWLDKxqCxcwfEC80pACnbWoSHdSD6idbd7BgGU4aXSaR2GjjKsRrqeogRQuMs9VLu
NstmtETalbX7Oq/PfpcjHpLdEWGgH0vF26aNIARvGPuB3Yq65cT85KripBS24C5euav3vRvPUSPr
FwTZ93mvvdVzXg72YLBaNBGN/BEfNyMxy3nG6avLN8ITbuNB9yJiEZigxSwV6UCPO+x/3wcFsmtr
CTtOklrvkNJlRvtQ3/tdaFpy4YbTp139z3sZ/viy0O5r0rJ0qWB2yM4SdVVPb9NU18/EC5uA6AYU
XKhoE18u67qKhNZsqezYzgyiBg5OWZdbJdNf2yX5HxogQvfb9ebeJMLgEMn3o5og2LaGKPFqEliE
6oadTc5Xw6mYAVAj7St/+Orw+liwdyATANVQZE/U8zRGzAOz2TvdgsY519M3vyKrP3hn8wyjc3d+
6smq6bVFtZVT36j5FdT7F3qFwPCUqiKUzckS7JQjYx1u9LIvUSGwdW5e6BH73A+EQ6oasFwS21Tz
8QOb0i5EogsAfvaJqvHuVvjwbbqVVJDEUM9+2symFSqSUBQ+zUk9bBPNnmTPAl8jC/1ajMN7qgvi
ntwf2JBZgphoVDG8TMRABvgtmutoB1MFMRuUj4Ldwpgi3Aug8C6iozVj6Viu4gbDTXzlrqgcy3yz
pnsMnVXIf0BHSAT9tZYiP9GtC7D3aXc3C/oOxigYpSJk9VQWEwu8PwfetJyerhZHHyUYghz4jemQ
ng+jpJUjfFO653i2RK8kZLCeIvhzcdkiPRAxUZ8ni2tOKeRbBTAiXJ+JYvVASVCBGd+Q7kiq6A6h
UanHQpYPNo4zDOT6klY81Q5PGnYbnnnco7ghl18XsdjmKFPnlTq8WHTari4fMIaeM2LttzV/K23O
O0DZT0M2O2SknVtMBcWkVvxG6UFP2Ej5YvZ+KicZdDWlQWGA1EI72albcQRCOg8vndE8IUOCo2Ad
/oJ3VvlkWEGuurVkdxuanwt8cQuNGOxy7WRfEjHsjQ+QTNOFacvyChpf9Lrw5V1Vx8VrZUMBwBkM
UwK81HvFLmGwFyjW3G5gLDao9YmEurtV6crCmm7EhvX9ul8s9cVUTB2FSWGdiPofh7A6ofA38sME
Cr/PiS209l8p0abdufSHhdsRxvhPLV8jmdjoIVDL2uqSI52mI+VOQB7eolF7ykUELemqVFyOc/sf
FdTL1mgxiYgAt7FfcqvzDXb3dyVbRdCIdKkOV5ozs1NfQ8z1faa62NdJ5A1fFKI18nUTBodPeOlq
zISt1WUa9bgXEvMa8mmecWBL2xtfsb29q+KAdPjgLUkxpjucd1VNC92I2dN+h69O9J4S+rXgy1Vg
poxAu2MNxxC8L5lMiWAWWh11qpLTN0wyun+7Yxt++qEAoKg+n35IfT4oKou3r/6Sk7h4iTR9voQX
5RnD/Lljk/njiOwfwlHfQCDq6xwkRJlKY1O8UmnEuo08IdAIK+zNqFGXLnpVaz/fk02SVMTnLi8r
ULhfg+fjoXZkSby32JNDzCnUD7RBzzlvAEZc/gL5C5tZ/f5s/B7w7FA+dio8AM5ch+KQUX5lugD4
o0o44edWWigu34eJCHOe9DicL8akGYVTKh4qeND9YjYpw8Xg0mnAkiXFv1TRrfAaCdJ98vWuAarK
XrJRg7Rlnc+9hWJZ3m8V1mRl3yE2cwI7yroOprueZTtkPeAQgKO3hkDVsFR3vZnV//o7uJFbwuTN
G4cKd2AOnf06gV91QIVg/ppU98d66MYf8bAKDyalGm6A3SYNB94zwmsDTqM8R1V7nqQmHpKM/aAq
xiwcT2YoyVx3378AQctVKbjqiu6uEZfKo2To1F4BXUi72xyCdoXzO1sKz5XiqYFCdLWiR7IG7EZr
fkbkLHemSqFWFcG5ezKETSgoNWqS2wk4fytgYzF4aq6WFRpn12iqJ+I7r4Ymp4/k50QvS495VfD/
+gN41O4Jl87mOWhOWAb4+KN7LyaNDN6ppKQo57xmMPxSLWLwDUw5K6jo3dCHFU4uLtUQzud283K7
MADfz7vwYxHJR+L+5dI0R03eN0TPIvsOWH+cuE/lUKkh3yR+vniF0NE3vBrTLL8kTygm4eZSyukU
ETDbDX5j4rvSKociBdIDdd3ofSSwMfuux2wBlkxDP3PIlhBp86lm8xLgHzJo6zADLrb8pALqgIup
4UTEQk0yMDk7EzwkpFyOAd9KAKBJD5LMAdpVmHHmLzrNyoRabymWwagk5dEoYr7ILUYYIx+i7KmT
+lqCG4bF4QMG+yP+BgIGe06+50GgHAleKJ+l1cqZIUNlXuGN8QrsRw8sqemXxtuosb0dzzIg2L+J
dpHoVuAR2Q+bzpQjc0zhNZsNw/zG8vp02+Opj+HXNGLvKO8mVQMgYj+iHrvx+nbBKATgHXiuXmye
u3FHekOggBZzTznn7qO2DIbWmRTS2LGsluVO4XjgVLT2iuG8MA1urWyDIYePHJpycBwZ2t06Cvmp
uqNEtC/u9w6taP5fzUHhCsFduw5dIZQrWpEVDL6/LBnRoBDEKTW3qKyohAI3fceFc0YKaBZipno0
sHmv5tTFwgBc54gC5vnU30nhV4Urp7IG6rt87COIn+/vDJPcpR5yiqJVX5aDqH6aNBcJLNwV8u4o
XdKZ7a4xX2cCq/KQQ1LlsEaMZgATZ1UBcz6ltxH6VKUMxhPeXV+Vf3qtFOlllMWrUZGIdjQvGzcS
7SUizA1mRqqHStTCGOtGJHBjLbkxkYDdYf+220TdIsYz+Mo9CHcTPxc1JcHkgkqLvFznqbRJI1UX
7enLXiD4ZcBRmECEbGGoioo+dlJg1ic6elqNbS6ozR9uKCINO5xhiiABDD3QYU+PXyyE2BpACZ2r
YvXcl9SV4KRFEYalj4TL3tWyJwL1GK+8lIEye7j6Nc+IIktulhzIQsieDrGY7+A3STaj+DLBjWxb
naaY367RUzczGonX1ZLe8Mj5hHUQgb+mF3oktrPOOnm4ya5qddWR4D3QJ5t/tjsucDNZOkMrURPQ
e2Ei16sz6S0fL+erSui8GYrDUbX2mFwog8fAIXnNZ1GRR1OLSF8Fdn8u9Oh4SVFtpmfhEUsBg2oU
HRADuOBtTjnBybRlZHzMRmx/E66PvKnn85dUTFjs2ZOwu+/NO02Uwxzo4E6DCbGwGJ7eMKHIzxD+
3zbbGWhsFB8LSJsE1Bc8YOsd4MhqYV7f9MrnXdXO8gRTJ3IGJt7oKNhCSo6kyVI/zLIMeeAIz11W
17sKbVGuebdPhDdWa34+53LO3nhYdvnSWIlVJdTvtYQMpV+q0Kon0dVQ04ynEIoh1RRKb4cdNT8H
cKdT9cVxGwSR7pFt0OOGk5pm25PpMKQuR+/cEFvgCK1firq1dPnI5rdkRMGom5nbtkPX8vm6bUOl
GnmZ7dNsHr8ZfGuWL+4K5IOZmuneqJZBpEIU/LRbI2gY3BOpKENHtseY+KyrZQQcZo3DQiUy7DlY
MQBYXaoQxUzP0dzglJmgdENxMOSXcewxolAOzVL2gOK7Io5ShEyX+HJohUcWfGJSXTGvgwoYMrHh
1odhCs6oPj4/fIOqXHsjKNlXneRFTHEV40GFuziXL/ayZqMWdDCMxfN5NV+IeJ83NdtwalQXSUHP
wLKWJ9kGYJ9zfkFHLDFikAF3RVd4qmt3MIZEQmILRfQqUxR8Y5wnEGFC2iR151vtV1ms9aCcJX/B
/GzYJfzSac4H64o8C+A0NGNsP7tWEB3IXKIDWXSzFdBWsR5gyi60AtfuUquvvr5EFD992gF/Z1xu
S1gNkttEjROX2MZwjFeu3eoLPPnL17O1INJF/ldozP1BVW4oxi+LEo2YSa5ierR3crzEeKp7elFI
1HG7BwQW0xjOIvp+N63lakr3m4gP/zbG1/8E/7jU5SZARpPC/99BUKfww0X+qNsPbPIF8w9IS+O5
io8IzAoPMZ3OhWQsu8OxUaqW4fWAMUy0MOI2rWhUanKC7iTPY+S+WYvCeIEGTr+CxEfHo3CUkNag
UQ157ZOCnnmOBIXE6Bf0fx9P+a6ED/UrA2eroq4VOC2uEb73bwpUwrDRRD88wd52YLnLEJYDlvtL
sTXI3PTe6cY6uAf0g57Yf3c5dkXBjt7YsXD2gfW6tRU6UYhe5QW7YMOp/o4rP4ii2HSHmoW3FUXo
ktvupj/H9PXOBA3kRP9qhAhLRXFuVDZsBRwApTpPTG6fkUB60HBgeDeVkaJqV4pVToZX8ndD7wPi
JSCVjJYRu2CEdDDwD1wbJJzfJfXxyyyAJA522tcF+gxSLTu6zRYoVNi6S4XUJbl6yEIymzG7D+pO
8LU70WMgswnBb76bxqX6rAS7qQZx1fG4slBL6+u0WpvBxFEh66r4WOAcY5Ku0Mr1IBL9CUiljuzA
AjdaLLvyluTl3IV35WjQE1OsKPQig9VD9YVVfD34d2Dx7ZdmtF445xxSPP+Bg6uKVMU8ZaST/lAE
3X8XQB9LQse0ao2obtRuuW2zb9NpJsNAXIOqf9GniwQnZRL1CfsAaI4F1e03+MIgoMHmR++ZMIBK
6mE76/AL8svLc7P2mv1Gq502843AOLnBcFC0jJ3jzMqj64Z2Mhjig8jUD/iKl2NcNch20DfQT9K/
Vebv5EK22e6lEoosoj1YpjkFtcDQJEcSONfNYj+Bf0kYVLnWqk5Z5bIed4vbrPWInI+nLrcXShxb
jgVcGwBzJyIkV+yF3A1hIuovDQQvMKXeQ+hFXB9m/beVdHQpWTJ0UUsls9sJp0OdsFXOnu1iKgrG
pjGODZOTS/PECJpS0A4BunEaeGBS6sjekk80oz37TDRLh549PWE/+YgKYT7fSgx57YxKxvng9X9m
nRU5u3eJ1M3iWRfImeFME04U7pKNqGJdX2CrSG0Bcw/asULX2Inv8kpNzsoZy4BQmruU0Sbnibfr
8d9TKFC345Xp698XJlGkYmazqOU6Mc141E3TeIT8u/HmETrIlZvYKVWfSjMfSNF931f/j0vKGtPX
e6JKnR+iSzogKGMqPwbJCDKShMAmgbBShi4P8WUszazdlMNgxOYbavziADHCYRIEin/7KfVUDZ+t
lJdZ/eLLpSPaaxzBmXfRAvto3ufUQfERrzTHYXopcGSwasZ77cHVHCHyEyR2oIjRMkwLEeQEjT3h
AZ5c2sx0bcv+HvQlMtb+RSPn7H2df6Da4KrIKKQHJ+aZipxcfn6k1VZ7qQwbGCHnjItVttKNkqCy
VXngPMnPcrIbx0Kf8ODVqZvFtLeSRRFoTeumGC5BH+y/6kmsvT5aF6WUFIJDL2HRhXDCKHPClkZm
KK/Dm1LDk7fE8WE484vPDXHRawcUxJasr75D7bL4Cn0UNcxAGYNUDG9DNDIFa8pryPj1+tPTrQkD
JSoJ1VLkxsAAcgr6fbcFC8C5onYY9aeq6aR1HSK+X9+XxVjzRX3sPGfM6WvQgBV64SoV7UADhSLM
mHoFmWMg7UNp6m8asuCA3YLAVdilkiqVYiKX9tOnzCSfaX3ele+W9U1pNw6Or2/3HAqoiNp5aHAV
DknVILAlkao1RVF5oSueGi30WqwXqcUCQAPFY5mAdyLoXBZITNQEcan5HwvkMbv3vTmlRdijwX5G
q0HaejuTNJKWOPM7XVc6YsQtaEKBkNhtC5tDzIYKwz4YXTB2wOAytSozCudTWrgQnBLExlpTU6In
HKFPCr1Mv79WWiQTu7mQxX3uG9U6rqAHJ9vCZ9Nu2q+ydK1ri1x0C3myU/5XyXs0a3dMVLjH1nFv
sDiLiDOhjtEQHWWK9N+sN94xbfgARPyJXwC8xV9p5W65DBbMP3cHyYGeBH7WvwMlweSQ1fvgwBiL
NCCY0wbHG6qkM/ouWX+0hMn3f3OJTksqiDh3DuuHET6S/Xdy31AjnYAKIqVvuE/vwFvxtUyEhS73
mZS4kApZK/dEIut0ylIZDFy4ZY/OmuIf+6N5mRJjq8P0TmOj4PEur1PGQ7lCgKPyo06aSI6wsJv4
31UrRZtK0sjVXsbni15yZ4fJMfzmQnaJkQpHOyvI8ChVjQZR2L5mwqgYKMkhdKMqSTTWS3biugYp
mCtRWx5Cj0jJ1J13AeVzqmturV7MOah8DqPApOlv3eKr6W3aD07wOKCLOPr6q37vco3R/Qvw9pdk
CjnnoCQk243oO2fJBQyk0X4bdDTqRuShkuVgQS9GoPiUqWHAqrzrS0wIn9/IrmGFEirWoUQ99akO
DyUI47Sw0X6At8zWczpQ1n3H/DWyvfniWNziz6/kpAxGj/I7cqGaEOJqdg4oMRqiuTMhK5JtWMlh
Hc0+IOuMqDjNLIwwJoofD3p2OII2n9Y5R9yhWESvwnMLEnSi8s8cz/Tl/MchExv+fMAaN7AnhMNh
hmS6qX8Tua7qUFJS4JR1305R12AoMGWrvN9kh5hxw5Cjj1KQXCa5LFfwtDcOSjov/96csK/pL5G3
EowQl1W2GqAEDNhYPcMDVVi9WtCmVsU+Xz8LBFgYnK+RpQWHTCzKfLVnzOcI8+3iFecmtNqla/s2
+/JZzjrlJsR+OcIJH8UOVhUwtV0Ds8Thcmqdm5f9+Gkh8ZA1N660lCNjIoEhLw2M1n6LAZ4FGS2I
zsYWDfGzS1iL7JqF3HrJkf+p1Zt19UDog2IQnFwYk3GAsNQky2sbnMy6jcwejLZAytyGjucypCb/
8K8Kq6/r3m02fys8nU9Lnma2DN7xI1ssHrxS9QH5klwdOIJvZ0Wtu+wdTkYpgykYukGsM1A1E6Su
0AoNr0OojBkiJeqqsZurwtJh+P9n3tQX+0qLP/DWnqh/4HGL/hXHv7Nq8u1fRuu5uxup06zxma0O
tSgbZUKCi8wE4MorMYXX3boGeydr44NftmOpwqF/lPW4bYGJgAdnDF5Z39meFWFOV4EBfX9RUh2N
ks62yaNjDLY7nv4spku4X+45jUj1MZMU1zbLmqzAMWkjj43QxmTSZgCl5Op/b7a4qr7buSYYQ11u
UyIhhXL0K84ghLpFng9EI/McehEWohnjqTutTn3Kj+kRBZMdvS+0NwpNSDf1dsVTIq5dwbbOa6wa
uNAHxEIYihdWn3vvxkDXzTo/e69QnPhwt3bLiy1fcXljjvh18HJGBuzTBQn0hewhysI+1AvRHy4k
Y1KogobMzWEZks7gI19zOSFZteSICLaXfeHBrPqYsBGYH/0VByTCiCwdkWx/flwEz/jjvXcj6FgY
nnzM3drt/HjnWTgLlbSadANtUqyOnVw1JQUemK3zTFfB00U2wshBYcrp6BjIhB2JjHhK/KaoLs0E
tnE584V2pVn382XtUvRit1wERZLRdJ2zH48vAzLmDmEfUVt8TZ8Hc5XaSg3G7gmnM2o+DvlAmOq5
z6iqP6Ybd09du1AhNUlvA0rDw867dX/T/CMtWoP5098uTZ1hbWH/FBhNpvw2/1LD3YrM7dq64ErP
M/0Iy3JN4wJVZi5XJLRA15XClzFJJ24bEG8c66nlcfLCeR0a3rMO5Mrv8qP6rpuBgPeF1WKN3gbh
aowOhzGiJGewSIKTKW10Oc/eqrAZCvfAfkBxtCtNuoY66FgQt0xwzXdFc4JiUwTb/zltGUG6qbPx
auevUe+yOluBZmDxnW4o2unpOqV7PHKSKdWtWVX2qRd4burdDWlTSjDbGWtKOLnj2YmFDox/VZVb
GYybPGp5HnHa0NkiWMI1GGukGzFOKhjhToP/IBweclXOChaUYxAct9QjuAmZrFr0l2gLhZDYuzfl
Uk1SQRj1t7GB0NdmtKCR8A6ApQNvRJCFpTQdmrr5zvfCNwIOZmTTLY9zlY0/RngmAZIdEQWd/NMX
CTOfCk4lvpTmYCJWa2DWMRxFz82Hg7Yjb8dY1NQBIQdUaaBf41YRIFiQ9S7l08JFE/OL7ROplcwE
kTIcQeKbppv//QEsyUuNORRRdzY2CxVVSnkKJ03Cwu2ybb6OK2SFl66jutZYtZvLUOKnAvIBbmMn
pwA1HuzB3LoSSsbWsoYOZ2zn2yM3T4iWf8dYYbOVfjo5bqzr9tght2lx4lbX0vti9Jecj8mk4ZVm
6o2w6S1a5J8Zl7q0hW07DPdpWIn6lR+LM1z/Es0T9+TJNS8GYPKM4SQ8dgVDr8bijMRn9pecQHNT
k3LIWvO7zOzLoKvkWjzA+9mZkdsJ+nqZQ2qnb/6/BuWSyfw7KRBH5Nsm7h5Q7wQvOo+cB0R32v4Z
1umIS5DNc/t8DGykirlfKkZsaqIHamTELNKF5oPDoe4DkL2v1eMiQptXCMhW92TP4WiCPuxMxK7b
ZZa+C/PlF+K3D1kxWmIV9v1ci0o2oF0ENhsrPRxkcwx2mtWHLNbU2oXGXl3A/+vsIN2KFGWsol+R
pkuS8WHrZIauD3KLi3srp5e6e+qgAk3j4yA289c91bbaLd/SmQ+ZxJc5XM3ik5QKfQ7oJprMYJxO
AVkKnrA2OYTqMgh0WlD/mi0rVyRl0ATBcU4vpaULf3rVT0AgTUzFpdFDVrR/wbpFm95DkQElJ9Cd
20LuIQKNLI3JD0gXA7GYaU27wx4EaAg9Pt0pxmGqBqIyWKM82U1FEey7dhRdJkDpO855B08D0Zli
kLLydDiSGygy6V1ZfIS4NCme2867CXlEks+HKIEc5MmJ2H67BBU9w1BjdWU0bEgyRACl8DKof/S7
WJ3IYzXtvcoEdyhVe2XF+IuifwYVixG/9E/KL+I4da9SsN9EsA+GZyDEHWsLxdz7hmruSBa7TRG3
bsrJUvsZZYsRONyofMvA1r7mx04R68x2j4Dq6zoe5WUEGviZ3+7mI36OtgZmBmmujBP8CuQNFetI
OL2hvj8eZnjOSlH+tpZNxq2Az0cPExX9YkAORhFuncMpXSQ5xqN2OiODqyWuf9IebHlUUG3R/+LE
NB0fLrVDJBk2f2bBGkbAkBKdbKhHXCVTD7ZONyyaHOBambtJSOwjLF95wTkHRZPct7Ag6+24fW5c
knOPGdNrqHksLVTiOlU2JanvF5XweW6SrfvBbTVVULw7A8GIS6UgZd+brZ2r8c9zwjTnrwG4bXHQ
BA8b77LGde97rGJ3rmqUq+aCkaCQK5IHWJP/6sPK7bS26SwPkxCzV+9LbaTNH3TkjUkvd7WwA3zQ
+NtzoRKx/sVJPZMkSJqbMOri+haFqiWlsWO4UXCfTk6QUaPjd8Htdsx2462vqVqDztmhSEMiOR6p
P7CZL5+RBEhdCAAEtUFig3lDN9xWCDg1uUOWQaOoibPq8N8BvGcA2Mx+bcz+KA4Lb/v/2PJbMWF2
stx+SICN+9vYpznfCThP/2wG1WQLD3IktXL8mHvsFebKm/1puaaxghMSF1DwQZ0O4DNoweVxA74E
DOns4A7ZX8PRj1hgDc7vSKYSF8O9SMnbQguPVlgQ41x91nrAvGsSG99253dRVS23wRyhJme5pHlw
TnYRuNMeTmcle7bc6jYtmJHDfF96tJH9hnByuFu9ZFtau2aY2c0qiFADfZt/21AjSajSlnqUuwrc
8exIOtQfimn9OIDCRKwwAx5SJuOstp9bwslZuXUxX85l8gGQ+P8JbrkpY48ueI+ndLSi64hxKN0T
9q60cuRZTpSeq2K89SHNEXWBsFNNNWRSBQDl79o7G5Q35O/qE6/KLdBSQbEGXC40XS6NMhDRkop8
EsBQD/Km87GtxFg8+ZzRuUqEHlHA/DRgu3G6mRDemyVRjopmA8W+2llRb+N8i8e8vFcb6ZQmLfJt
N8jZjRInZWrki4jymoM6v32N7LcU4GwdnzBJvPLM+AlM++/nM80Zlfm81BLheoN0j/JC2nik0uwk
r5LOIx4fBVtqsO7QitZKd2e4xQwN2IDLZtN7/+FPY824tKS/XEvliHFaubLIZRJu2es/tMfmm4Ht
7f2euJ1BGxcVzst4QdbGdyH1qtJSg31YJAc6W1jZI8snl7ClWSj6REX1KtHxfTmiYPenXXiGJBrq
uM/OwVsNqEZO/zYY/u5hD1SS6pcoBWDk2ZxW7pqx9IwiFlq+vNmY2sDf7cQwEpNdKv8gGaeD8iiQ
A/aKnxhInaMITRGcxD5ykTYwMvlvOwz0a+HfuMWrJDOONaU/nF9z1mIY5L3m/a7M87OvSO17Uwan
FscyygH4OfZTFsTbt2u21MWDYf5aNHNXe1ZikI9iy5IyXHonf0+Y8uw5+Z5VbAyc93ThHmhfnFOY
p8mSh2tOypymrpmiNjSFNbOOx/iIuObOBAoQ8DHvpemUNVJLuJ/ZpAMzxUJsgsULbWClkQhzocy1
wKIwp8dymfciuyvDb8pHh3PSnoX79XQM758nzNeNUoEw1IVB8TUwbySdd+yZ4DU1Q8gpda+YO190
6bDQWRSzHlOfG42nfofWUWtjSfodggAnAzuLMcL9/nZKIzQKCfP47cCKrjIg34EQ8+MdGoUfHIVk
uK9qW8c4mDAZk5opkJ3DWeltCXVS69DaZmfQX/creF/f3VmRVa4zYurN8tvjgGHcNyHCfefqYKNV
N/qDxbCY9rHsLpCeNoa/7g7wcwhHvZxVF5bvDUHW2lnV+tNVtk2odv7NiMXpr2LYee8ayrW2wDn3
rbFhKs5gv/BR5k15tfoP+ReymJkduL5fRDdZSStiXL8OpKm8QDIHbsBbYedoosK2SHfXcQ1t6xfc
hz2aovo95VzKhqMY9FbKk6wwMrZDtBsqn7k0z+BuaiZ/XlWLNs6jcbZMtWJ2cvAEDwdlYxfhIpYO
OEGUuZMjDyrodfGiAzaOFQ5qHXg711DU5m+t7F5eqL90WrWxDrbUfAfesIfIhj97Gf/gtFQhQ1Du
7uHGZSI4dM8fBaa9w1YA11wpF4TlobPz5UcxeNtb7l0k8w1fYc+khO6tk3XofUgDK3HqXVdk3grt
p+/SeNbsLJMzVj3gD++mXUWU5HvKyfyoq74kQp7jEgu75AD+kCU38SHsUEUIcarFwBsekGhBAofC
8FA8JUbtGLahePofY5P+LtFTAIK70t2BWHUR9PRS6n2bq88l4xYduy1flxJTPdgpyzYegjpIef3s
AG89COVLDjZOz/zk+zATQI8hs9h+ccNDiD2LyDX4j/y2NXF6ADZ4WUAVSCgWSi48FpXmbQjtHle6
IcnNJ0Y/pJEmJVgaGBXGxgzXgRX30upndwHxe5fTx3PLb6HBtWvGhsF55y+p2mZTXXvA5u6X9j/6
BeMqJW0WLsrMRb9tYL4hBaFF8LFsCVR/iJy/PNle12Ynsva3vXnIuDBs/0eWUh98YfzhcVdwpuu0
dq+TDeVg0ES/CUI1w8T0fDHNOyJ+e2PmMWXnRFkAtNgQo9yJIcKGeq/je3d8X16jECX7CYkM3y0q
4BEKGme7cySxSWcccETExG0FsodQEGQB3ddIaH820XP7U3rTH8WFzLIaoLIbWjAtuPBmQzTMGmIu
PmvoaCLVSmGhQvsD22w6DAJ6z2ciqqJaV7M5lv/goGexWZ0zF+2WwXgY44cXapKy6tpaQ7gbUTDv
OqkOcpjkKtY1OPVq1YE9Iun0ZAaYVhdfSm5t55pf6+KHxL4oWg9+F3DaWZVgx8feU/dEK2QhCwDT
7ZecnA3Q0up9+AWdLdB3sred6d0Wj97jAEmVi1OUtCRhmwtui/R0k3TXi2vT7bi2k9j0V5JN+4kE
8ke4nPa15qCCYP1wDH9I05r1ZOqxz0OapzTzX9lXYEB4NWFA/iALJeMsfpDk+hDgPnBpYlYl6G21
be2lYh7TAEqbrK1o8Bc7e+Yk+NQwkEt4BmXAfSQWCihSXpNtD7aXMWlANdl14HjJpDgVIv/5xse4
5UxkjjPjoFnPC+VqeZTgJZYWSKAAh3Csu56XSB7qFy3AmfK1Hu+dkY7P7x0SYOIpBuIpAdhmrTAO
/xwdTYUSyfynwsEzfQRbNnZX/GuI2pm5u9gfQlGY0wNxCUkbtruBShbPDz1+Hb1xCcR+unxAF6q6
oxN5K3szyI7TsJXtzLidqQDoce1/JxUZkkaoQ+YouwLH6SI/rJz6Vx9bOMNDEJEnFGGKnVhlIUTY
vTcgOgBtPOeYx4UBMyrDOSqOdK/iekQL56GvkdVBIMEfexgpxhzZv9u9/Wfmi3+fm9H5rTObrzAi
Ndioh3C8NfXbniQddmzi2UBggBY0SsgA8aEH5v6SzaLNGe5yUI8U12ZwBtW6ACkyfQ+fPJpYvpIn
9UhJU/rxKWMNOZ5L+gBSZLwx3yB0R7y/1nNJnG/0V9KICh7pTzLVKT03+8ZVF3KEB8qa7Nwt0BZs
lLDglUYXgIZzfGPPH6ED7trHbULpHm8jCch4D0hz13JZvJ+hEtki00z7F3XH0iEWlUIXAp3hnigI
R1Zis9i6MLHbXaVimPMEvmpaqmTACdh4hXBHY9kZVWXP75ld7ZYOBP76dpt+TmPSuTTPk796NKdk
6jeBUENMcHn3RZ5+odsm3SiWK9tSoWpF1qtvei97awypWidHpxOK5Fry1CL1Q1eUQ4RO7ertHJuH
WuYAaEwlPjlTdwk97hPxnuAmVywe0hJQUk1cUC0Pbb+8ei799Cqjhp221kfEgVarcb0V8a37MepP
qUnw8A7Ka2DTVNtrpJpZokIGwvK40wIyQaf7km2o7OT6kpF0sZ+g5uXhEf51W/PY2hj7Y6q9HHil
eImgTwP7DVC78conIT4HPxjh45gjewlo1+THHPAc1DzdKlF8mIliSKvRJalunHwgOrSJueXE6EF9
V6/GSwgnzM25czBatdRVjgjaZmWcy7vRKP1HN1HLrzuNokMEYAnoJLEnqLItoZonJPmoJv8rZYjT
LAyOGC9SSl1EiNX6A7c6/3CgMEngoaxW+9WsgpOnF//ENwUNYv3u8cnIi5xE+ygE7nRMCG6RLIao
XMRL6OR78sizkzEv35vwUTEcCRmj7vwgTgfcI2kLZeUWjUExdzVxrR423Iy60o8ws0QActzed9gM
Jrjii+0e2yH490kPN0ZBj3wYZmB1RUnWMuecKJuhZqvEMRRezioLvNvxTw3Cgtd6krVRqVmFKHTi
VqwQYAomEZ2YY2LwNCW4KkLArQa+A9IEYXU83Rbc5QIaiJyXFLNSGJuLJNXxg4e6har1izZWVGFZ
xfb6g+cZFAYSc78g++jyqqS2Idfgqr5CawewzgqD0zia4i7kMkXEiblnVvzGcv8FIowPSfTDpdVC
4ez3gCCFnVo1I2/Oa1CxJdbWNTnWbp+uU/jMh+544dUhR3V0AZquNxdVw+F2um2USOG/Sj5LG6MS
53RJRk/MaTR7laXGhhMUFVYJoldMMeDFdtG3wyeaFPYpoa5QIwv/fvoS7w6V9z0+IocrQXi1vAHU
uVPV3DodpM+MbFdLcN4fLPmeLNR/VZ0Gy/4lgio5RSQ7d8Nzz909ok4+uV45z+nvWa/4oQnUsYuN
HgCJHLZgo1ydf4rG/WDMjVduRpFjGwTCYuQfdc0pIXBB+OJ91iyaPIeMZAYXznUXwtjo0dOrxnS0
NFRSygUVJyTXzdNfh15WjhT+I1fbAwRYmLRFoFj+aqdTrI89I3+evt5xYcLfofcvW1Fvntndhm8q
LCPhoRgFAXffamOqriEQCUXbq03V3eYwlAzwmWhGHUoKXqbgyx9Z0SFxIIIV6fkVAnNUjP+7FZH7
+33qeq/xqgtA7Htk2noSt8BubbohCU4OF4ucEpiVudSEPcFoK/kjvDbxgcdPZL01rEOqJ4QKhOPO
/JAWWPIwcL28BaPgit4eCn39nGf2MrOXE3Dzs/C7roAePMPiIe6j8yOnl1W9hTPx4bmq120tjCcE
dZdc+2z+hSvmguHocxFHRMe1IwDvDqv+rJ4oZuAOvKVFYp5M9Bb5EZaymvebIOUGmmvQ8Vpt5LG7
/yQjXEpdIiS5rkOiA7CrC0z9aOtr2nLSlu/RINqetXBedI2DwHkSOJ5AwZ9tUKtx1uEZpN9aSiRh
FCofI4rcbdQs44CK4nbMXg4VKD9yH24CY07OicUMZAp9VUPsRcn7hBJj93oS4hlinjjPBSPGH9Po
ADIJAkUa2qY7yhAJ9cr+eKfIf1jCA53UrojGodfRg3huFhRnNuw4hl7d7nWMQvFyCIgAwhpOmI2E
8rPHgfY8W05ikO6dW64zaFLpxEcY/uNM83RMhjppmZzVFlwFmZAnkJYxy2WxRmP1eGXCJOx9cLPj
BQJVh6yaLNac99ScG/BhFnCfaVjOIGi4XlduUxwxnBx592Dr5X9+mMilae1a16AtC4SozSqHkOkS
qsbLqPxNQJT23+Mz+2oA+OcN3s39AqwB3u3bQRzhbTH/Dd1AGye7XmHv4lMnr7cqFmnHmQ04YbPW
BYY3E0Y9WZLSskgOVwf3fZgQx4IaJ+qv6yPzmoiPh20Gb3yk2ovbSo6+twCXGStMDJTYR4aLzNxK
Wy+v3toAzoBydumy/wHilNnv/rzNLMy4kBRMerBJaxQVV8E5n060qgQBeB/eG7hGMAH3ng/it/gA
RGTX2RAoFTwqY/3grEixP/DIv5cnsQcnUDRNL2+mUb3DRxWyXUS+0OAHaEjBOxnB2w6MFMG6DAfN
vIfi85uhM9DiQowcfjR3nQ3VsDZRh8Ag1nTSY7PEPwZdP8bSlkrbUm+iZArtpayR46KmPYPdNS7Z
DgfP7lnLhpH3yCxMXmBcl22LK2UvwYn3/5W7E8L4KNlEu/Z4Ae03BtIivTqZtoA1WDH4lVNyjuJH
Xrvq6cECe4wyw+ChYI4Jcp3A/CybcZOxe1eAY44XSQzQHqIgB6doEndMrKK+K1pcg2BZrqbxFBmw
C/ESEA23rwslZ2KwpOibS70ZjKjCmKuiuSqwEthasVOtNKLRlXIgtyC3Dvk0LhHhzWXHD3V7W7xz
SGVd3KCDG4KNyIIUF4Itc2hHUX+dtFc/ip/i2D5XkPNtj2Y1+Wz4zA0NkE3/Ndm5PsgWMzTs8uPn
/2AgWJZycIXBg99MvoMZc8QDcMARPJBUwCJdWBMnaLvia0I7U4/Au9B5U3h4sTGRTgJ522mJJNUc
HpQaoWYTlC7MheLSGEbDjMLbx5Y4z2nws2jyyWJ8b4yLEgMYQ2EmwYhPmQSTUiTAcuCi8+oEpSnY
z3F1rTkgHoY+aSrIClvL3o72U2AfpcgJmldIh7WrwR6J2ZvIyD91ML4rZBeACId3op+tz5QKN7VZ
qzhNdLIBRwOeXVYVLekI993GkRMJkloLt7Jj3XsGoUC+gAdmzODl0x/DXesDOCKaMX6cm4rQtVa9
h2Znxigb+hBZHGYEFUCtF05424LbG7Lja4LOKJ/tKUylwwzDGwNFXuDdcw7yPxh+6HNHo2Zngkox
VEMO/dollyMuFJB9JX4nsG7NHM1YzdvIu7a6JKC9Kdf3cydch9ih4X9N6+EUL6xy6pPiRpYJH0aI
Vh2IMPOsuQdAp7fA1cizeH6MsAnULirloE3h9kwMMtFrMnE300kg/dRCzjNyCAlvvE/idq6wYuhe
xY+DHLUtjfhLJ0S/0qI4fatkfTsih4IOGRmpHZQmKb3cvLT45eTUABCv5pmagfd75AbbU1ozEHXr
S49yVf24PVN6fipoiMv6V8HrN8WcI5gsLBy5U9doG+MAg0K0NAPwtusjv4yojrDzAONaVaA0LdDr
AhJ9owAQJQ/n/DfpSB6ZCDlYLdFclFo1vYy6man3wEI/1Uc7EawxKKivnx9IatGlbEPj35pfL4ZR
1PfUBHBJ7EJS/nuRje9yNHUmnHoW2FgmfQdAnVk2mlBaU/qmCExKdobEtrU5IXz7yRxu1fRT7C0j
EKyHEI9Qmio8HEeU6OCp1Wdnr9UI8eSHN33myNMIR19aAkVCzUGTR27qGJpLixBQwwl8HkKT/LoA
vbEGO/ge7GrQO2wm4Y/aX3loovIb5v+sENnzZwnop9xHoj6d62h9bArjVdqqTOvsNuyeiq55ClXJ
FMpioVGTMl7AwIKvV8oSej24h0wFJ1wbheDjycf2yE4HoXGk2rfEjR7N3epWtmT4JA+x+CgkqGiK
/LF+J82JbPDVKskXbsgnvF2ofOQ1PRA519wJ+vcVreGoRTFWJ2HP76EbIY/KnfEvcoJSCHRLN/sP
uNXmQv60S9A6zYTYgbJP/IKuPpdNkFOtQ+dz049xMVAvf/UbhHGZBtier5WqvMeaLQfSL+YvtJUo
fmB+GjN7ZhPSXj5q/S+sz/6NS+onctzmYaf+NhpE93V1/R07a3fcxGH+GhPl6VrQ86kWTkASSbPQ
XZPVdZzO8jhZdHlxtQBo+wFJFiZHYluUkm6I8BMnQmfR1LglbD1Zh24osuxGROQYBk3anvHfS7qj
27i2GVXKAXDok002JJLDcESlSVvkYIHnPLbLyA+M1E/wTQpCANcjl1MmfgjZJ5yerJ/c2JQ7AUMT
+VC4XWDhZXpogYeVJNiHZrAxRoy1TY6vSgEWmCpmejNl/XNzZiTOXN3P7Lmg0NlNvtnLggLlvsl4
3KFLE3arY8h5tWNEkaBjM63K79cdXAMhN1pLKrMT0qRxHEqWOtyH4CraUH59Ok0QJo3n1MtK5ZeZ
1Ifql0Xj2m3pFhHhuQzsykEiRQG4LRdqrWye+zrnSl6l7Hh/h1ae6fcFL+U/ietSIkVC6fHIBA1c
DyXZEntJlsscqamGjMEoWqbmGFkxhwjo/sQrFtRoyn+Jxd/Mm38CSEoExXRM5DqUtX/izRjI215H
W1OhN6rP84C8BMr9C2Q7pqWMUVZRqcRsu+mNe1Yl6JxVopACA9GSsop0tVWFX3aWLrtUnQbQGtdt
m8xfZK/Kkm33FUWyxaHcQ4qsz6n3nJ/SK9u+vqg1L0agE4OgkhA5puOJkaLAsxqLLpC9a+xudwib
Vm7/4UXaKj0yXFSXL9EZKYr71EDqP1FkGfeovVh2DxNy1Xr5aewO2IoWS7lnRN+Zvv8HgHx+07Y0
IwWfXnjN0Xht5arXsmNfcaTSIZ6VohSOqWIv3p4+1n2mha208uoMR2VxZlyfcgWJOyuJx2+z2mev
xYnv2Ii8DR73ROJkWLvE7rHIH3080jeAUsv5F50d5aGJqBKr6NvJ+T9XBrSYQUqXrB38b029kTzr
aVlM4VAZ/NjzYLDnuUVSg5kLz+I6/F+U+Yh540LqF3je56SOhgHkA3XYFxO72NpuleGW2kBoN3a8
rz6us/LftD4Q+/zNH+g+mRrRNXzKWNAP3TpyCEejPb8BId3OkOll1HyyEHxHs8VKYzYEC6yVfy9o
u5AXtlau018pLnCBFCJ3Gtt9Wy5LtAT3W1zb/EA9Q35+fWo7YQRg8g+Z11sWiTBgbG/pMJnaLAMv
pBOU6b/WEhogET5qJkaIRK18zYMaZ/CS6I7ExzfFX+gdB5VAuTMJPVbSL/h9stoa22LuuQtSYbko
nZ1PkX+PvHbpQPizz7X1uhHkbfs2P5Iz2nLLihihIynXLbh/tSwt1GmqiqjHuTCW1vqxqUfGaDfF
6EpT1Rj/dlSH5cRrpFwIQUaVZ3vlhnwAMaz1Vm2aG1IN40uVhOCBm5uTrHxOHsV5QfflUapHZLth
ZfRsbzvBP6BohbiafhyxxmSnr1GrVlAgH7t95Xo6WIQNeZq5KiIIHZrjG2+xfjf9nP4zR0q9V/M4
czHAnkBSpIu0c91fmFsr+5O+MaWd2UFeGU3D9+ClMWUuej4T/H+Kp8hcZypudP2WhrtIU4eqnjQt
uJgltr2d6LsKFs7N3MkrNZ8QzWvJSFQfojOYLf1xf70qvMmXxHf/BAvQbZTufgOHa4dUPpDwcyrN
4aY3J7315P+soqDnDR+VNwuvpZIlqlxZjFWIjr/VanDyoZBlurFN029G5ecXUalPXkmH7eKsyLfU
L5KOtN7GaTdQWG2Xdasmixp3hHUxwAfvwCy56HK3mV8Lc1FdG4NGz8RSFhq/97p9iVkA0YsrCJBu
UHplP1keNFN6vEYhpwrQMg9cgyV1MWikeOnzDLWj63Owp6wR2krK5wKqzNh/yGH6xqnJ+fUvJi7C
ju42tS0HYBhdLa0LIDiY93aTvXB9P1ulKK7+eU10jNbXkAcjZlb1Z/5vjBmUSuhC5npEmX16rXzO
7vqaAiKkDlrzhATtUlVkTuclEsSDiawVXjrVQkwQmDPobILqMFbCsoYiHRpd+s0HdAop6V8m8JIv
bvw2KMi9De+VnnWZbH3aTHBFYmE7ziV/5pIjN51T+PVakqTMLbeHke/ZUTGcyhux9glM+0C34SG2
32Ui2v2Pf1OL4985qzZ1CWiOZ48e6melz6dsB9o9zKsTeA58/QiWP8bMHIcQkkByqY2TAJnD6+cK
lGool5Jv67q6jLiQJJ6A8cXpj/2fipmvNtvcbnR0vf63htd9BQlVXXB+It4oCWhTRLgeqhUqM1Nw
fFI3YLZ0aclunSyIw12MdqBDTYtKlBYz/0q+3iNWYP3//Ag6uaxfqSzpXQkSfrfH8+dJ+SCJ0WQg
5ZNQUXOOog1nIDRyxhoZuXY8x46rauZ7YAydh/Fp/kjIqck3DwTgykz2IwaQflHTaZuh6PYHYOTi
FRdSW4KGm8mhpJc+FsMw2o62WFLWevSxUWuoM2XbXBYzcmkmQSwGx2YV4rJSd6xZb1HDr29u10bj
UwEu4sch5NgKouzye9ta+YdGIxuho7AjXFZqedlzXr+s59pe0gQAWLy9vf6V83eT2nW7tlNb4CZU
qPrUCYXD3ZuB/z6p4mWeT5QIbWAvCuFkoBNTJfdSPKjSpGwn5NU6zjmT8hK60CcP3aoSnCuvVBBt
qQCAfPOarnPGY9ZrfRGVrP8jeP1UMeJJdWB389G4rPslUExzRrEq5yZUMLKz0vPkz00L5jf8uD2G
x8IXf5IRZe7+gRljcBPmVybmiNmJGtQmh+z3msP4PLHbx9K+sSaJO4t81vn9z13STgG39fmRPxon
BysDdbr0+zyot4QQNHTVV1NMNldcQ1mzLmMRgZtXM1vQOYi42EqH5vZK4bqSu/8mui2cb0SVo5os
X7kP7lo/S4hGkFOadz9XQNuriE3whIG7Wa7R2DF5JnAou01y4AnXRkBkw3qW0JRXVG4n8UL2vOm9
wvrQnufly9ZPQV/fLNiLF4CqfO6igcAamZrMuErWjrvkfQjivjK2hLV/rm/iKiST2dxWtSqQgrKn
XaaSYmMhNLW4R7mjRRg6YQxVyzEu3Uk4YvwgYpmuQAnxlmNcMPQsyed0dVlG9W/qFkKDiYgC7egA
7yPzTXBnDWZDbA7o8FMK2pM0NvP2llkp5F8eKWy1SBAJwWH7n30q1uKZKohcUMeeU7z/WYTEHW0S
WcJjO0sbAh5a/9GsTse+9Ln0HNvEbjfiV+R8aoylhMqlle+cFtwYxYMNiY0jgoUwi02rJKYL+Z/m
b7ZtktvXYZf8l+yswzI7Jko8vmGE8nWWQAclLj/jmJudt7MuTLqmsSwv7LcyCnFspBqPOddiX3As
vrxnUiAmHpxJHn0tcHutrwZA9dAXBc62s9ydUd2G741GHg8YMkyOWDQqPUk7xsuo19aoVuf085ft
UC0apQItG486oIMlEOAVQx6EcY8OZSbWhw38BiRjtq1VE25ecJrskjKum9OFlQqEPsSSkcFjIC0J
jrgGLvjWfNAZBadCvb/S4tg6Gw0TNOn8YAEk7NP45S8Zqe7nL4oiP2a9q8vJestN5xfqfd6SSw0I
YwUZGQ6c9lAkkbq7pwXMoeGoI3Qi+Tr21lQV5jaHLo15SDOJLN52DMBi9IKHflMZ3NL9SE6e3EHo
GK00MPn/V8Jur0TH1vw17d+S0h6m8A9A24K509j5jeUM5L3Y3z9NaBYmP8RNpYjMeuhKXUwkmXcP
+F4pgjI43D6eMat7QVa7MrEVgFZAZM1AbO9XURMEqi9/HaM0q/Nwy/xSzdgexSv555bafTobTlFd
kS6GxRZgi7IWkkzijDOwGZZ2qbIN+mJQrR6I0ZVYAjNe+8C/5DqhsnT3s9084A/6c7ZT8KJcvkjE
pnmY7gQ1MgYyjPQJStfrHPZLKCqKC9iwozmIUhTdXMnZso4WQ2wvQdn6GfL7Uw7FXKchHk70Y4n9
ZMls8d3HaZ4x0E+Rxnzg214SadyB7qHhFGXJihj+QZR5GEfDCtdaz4r6BBY95OpY9sfpvnRZKsNj
ougQokg4GHcjYlwCk9k+rY9k45IITyD5ZTvCw82gtngYgEZlMwdoEQys5wVmyyAfzkJBGSb42ViG
HTHyTZbdodknpDqOr1abFTUyAMRH4ppyUZF0g/1dQs1CZBITFbbGdn9HhqkIIxkONzHxu54Z/F8K
9gX07J3kU8e7wYz8POQAOWcjk77zRba6MR+DTt5wNgqFQbWFljsYa5K612TqDmU3ZpIofgjLuvom
Sn1s0+aQC07MELO95Se0oEAOnAKvKgqIupR1lFqaKqvm83pCqFf1n6qsLAs0h6zlBwbyHXUzJ4qR
k1GMVMfmeNNKerXLdC4s6kqCXOFkfDBIcw54l2YFry9PNvDEFwfaRarGcB35VlAAV0ZyRXl7voPH
VdEJH8U7ZlfvShLfgmlTj7pi4enqzeSyHiJoNyFy8JYKGUNAAzIxAeoJv419pas+sPYFJQ5uJZ8s
FXslR1MQI66Tdi2H7pxmP6FRGovkPT11LCKSUIdubXLc2UEM4GKhzmaF3LQE/R3effLEAMpebulc
1pEQjiSi86iMZkqzkFBj75vLVIzH2vY9QNbwfenMnG/KzRDQq62Rl2uWlgo9n0C+WhxN0HP5ZXAG
P2j5q/SIwZ0QED4dnSP0SY/qC8I1+VHgsMeRC6DsmpwNjtdfg7IznsonAVeXm8C9u6fJnEbPg3VP
VqPWRTzSbsB/Y8gPUUxNULTJbBesSugHhy8LHlvSLBAKl1Ksx/J6vC9znF+no7itPRecF2fDuB20
GxotD+6IrBhTspTm/B6qEAQGy47O8EAqs952q5icWr3NowYae95nLsASzp0z/Wbyr1CJI0qoYecp
sGYCcuRByyJYV8HwnFzA3ymrpvreo48fcbeSjdK4ue9Joy+bPTsfQ96Jnm4mbyJPtemNievvYvQ3
LfKG8ez2bm8tfLDSNjUWVkl3FmIca+AqspaoVbGQJrF68PsoxJL0ellxzxgEUZ/1VndW+Pcr/Law
TpOgR6WfhIVuTQP23vxfc/SGO5rjLJ7/Og7EP55aif+iDFVInKT09XYRHz9T42xeGJq0rZc2E4z2
wDVcrQ9EhM9BNRBfUc9C1OScFyVPyxVH7BUmxryKdnWNNyKQyHQ+CT0dB3m4kieLq3qLj54VtZvO
dWlyWcotdBNBeyTJQPwz3W9EvnostFiktEMW1u6AHUknMqR5pDepumd24zx9xGtF4F54tycFYbXI
8D/NbK0qFeulipfmU1r/uv83SuA310yCqPX41XoSUugHEsNPQNGFYQ3FPURCXBda1jWYQ5cyXZAu
52aNx3AoWOdyzpdF+ErYNuBTVxukw8QAJ2cJjGAGeR7mNhqaM/rfzxUpw7vDigIlofXhqp6I7fAU
kJChQm9V/exLVBTMamDUvC6wSAMwazJBojIWtK5QlZWUBJpq3Q5fh+mUnH5aQj3Mff76ASGTPEx5
N7zO7LoxhXZiJukxmTdbbuIAkbDiQhqHyiiuuc4VPQZESF88w5Y1hbKm8xxZXZsGahitaT3aV3VA
A7DFxza1RFtkdoWn35FVSflUVI57xdgFfhbLrAo+MRmKFCW0eIZ4IkLMLPtoo4hNJaTBjxBMNxav
Z4ZIefIvOxR6sqtzp7RH3Jwsn2VN3Mr8PSKEWoi3nRUfVpuqtZlEdLv4JaW7f+SydC4H8FvsD8FF
Rm26BC11k7foQWiYg8LDwzpCusaMiYplDH3ggdmxVh+ZMPt1jn5dsoMZxCENovfD1Lp/YbxCJSp8
b+dxtFqJDm7VBhAPCso71dIH+Owitr7Kka0Lg0d9VQciyFlo1ohyaD6KEEJXFQmqqDg5r8KjwVlS
yU8STaLN5llxwkeGcfyEy01ZG4Eykr6dJEzwyUGxFZTDy1M72dbSARczYAQVFNsY3tqe242ytjrm
Aem9nYuv6QocJiLbiNhOW91fcEM7DlHoa03U/R1c9qmbzR+JnMnmQLeSmGJKwF4fr8s0uEfHLoR3
wxVFViOMv+euhb0i2Suv55vtnVf+u26vbkapKPd/EjVpLgo/wCYTnOgOcA0W6JsrDMgZoNqyRHVZ
KwoqLMbpe3tjpxecUI5AzFnPFmQZzRlOh5uW/RuMpx3I2jXVwjethG8pSpjDafCaQZBZXlf9SMhL
3SWMsPLyecjhPo/dPGGDdNRZiiV/YjACC6un/Wx7BwHgnsshjdRwRoYe8V5tPsT/xOSu/bFU/lnr
QONc+MouMuoM0uoO6NAjM6jL6uCO2VuI1Nd19MRtudZFtrfJWWqzZv28wvl0BrE4rYfdLMb3YsmB
NVyfIR37kbyYKvbZJdmjJ3ROR8JY49N+dNTB8ta0v1FQNEB0MBUqyEyHteH7U4lyEJpSG3FOCjJn
YsJSarLb4CK56v9FlYvWp69tx3KN/Ye+bEeps+2cRO6QPTqtodSKMjpIJAAhdsDJvOhUT/Ys3JuH
0o59qRtbq4g8AIUY4+iKo5PUfUEt5lLtLpqJHVKmX7qG0ZxZ8AeoKZla5Xkm7MYI4oI/EIYjz36N
euSgwPgWw3ZWskINsCZoDbw3VIT3qU3qQa487vQyJAK5eh6ljHTfRAeSZNqEjEohEchafsPO+Aip
9eOHcSaFrrjhC+yUHR9ck4Q4yKz0lc3PlqJvbRB66jJnt/DIrxdEmWYd7vkSXe+/nTDcSWVcHvcU
eeZeeRMSL6ErKICnS1Bdkr9aENrLZxqhOSwpnaFsFzsRIM4/lwVVIp4FmwcoNjik7D9y3Q2RIpsc
xd5u2wyKD7Eqfp8yZy+/vLuiftuw8adQwlX4M1RqbEqn4KTgZ6SXqHz7IB/pi8CjYa5LDMXe5MWG
ulsVXyHcw5w2Uc2AfiwHy5ltgkgcDv6euF9c7kEZIYeOZHxUK8AOWQsqgonE+UvP8QyB3mqBd9cm
ZN84bEpguoX94kghjhfkogWxICOkWwrtQ4Tet0ChIrFrGre5kIpdw1rTt2Jkt7R81e2J/KZFf6BW
RHdbdP31u5jk8NjUyrEswv6d+fgtm/nmbHQBEU2aWdIpReKxLJIROI4LjBfNwlnJDrNZZxiiaHO5
091NRwcB53rjSzY2pM5EOp3NgBo76AUVBn77dOOI51CVqlpbaJajHu+VLWp2APdSWq9olBe77wBZ
29RJvvJ0wQuBr0cZrvsk5luvqUiDqoYemwZfqnuKGbAeJ4lTiDN9Mmh0mhOF0GUG8KPoLvSSgsIG
FCtKQ5rFJrdU8FK8udJjiRFC6G7SdgdfHuxdBLlr82MzlCYGjrpnNNnZU6bc0N7UqmlEWBG4zpsl
1qokAtswA55J+Ls0vwc0grclK+XLNC4xip5pRc0D6wShblxtrq8PrzL/5AVHkbMmKbBpeyAIrtBf
0CmKDlVvHNalsHlRScTcCUZ2izuVDLC+YeUCE1MWfNJeC1PQv9FfZIjs/sLM1Wy2YhwVggmBfmLt
nDgtdxnjycus81p20fQojlw7SlRlcrQYM8st2SaNj8zuRg7aarZYcpcHBABUV+adOYxh5evYXbT1
jmZlo2JP+JpGp+xsz/HliLx38eNYjso2PtdyYOIi/bInf0ngpaS9ual7lN2FedxeWVTLiKeg1MG0
nioIS5VVp8b5ydt8xAn6jQJsCAr69TpRvEKzFE4pKJ/micBrev6bI+5yV5PJAd+hP+Dw8l1qZ5d9
H7XHZyanXZzavNtzb63WOJmWIkkRMt4tjQEAK0nxrpWkjKITuArGJ5DS1PJIHV1BHstIYdyLx4Yq
w7KsuKOLrVYhc/lK4BH+vRx3DPF1FZH5DZeeN9P+XAo1BNB1alPTWHbE1/Fb3W2btPYxlAx7YDpn
Xt6oec0fY3CRU/qU9cqkJz26SSOw76Gv7EkhO8KCAt8HrEli9NUpoHorGPfuYU0ypV8Ss0pIoh+9
0Xz9mTYqd0Im3ar7yRJaHXImSZR1f06GZ1mlqmtti3d7mOSVvD1yBgRUpz3VPVBV3Y7fBcmhI+1O
eyLcH3LLxxhDgvWfInHylxReyNVUxPe5y3DmukSAnFSs2leMTmMcy6BCJZTF6SF9HOKT250v/f37
qSPT4rbFL7uGba9mZS7yrIkyWfjTlOx+BppMzN++2r5RsxT6sKObb9ZArE2rC7vYcZHJiG2zei7m
dXlyYBeGxxKtx3whXT7U1SrI7Z8i62hKT5nX0gGrmIk8UOAKdUWXZtWi3C+WRQ3nikviJOlg8TT2
6EbsBbFUydU86yWXOxZRzZvBz0ah+vby7EwjKCzx0UCZz+Sc5ToBwpXRJGTTpvOnkJ2c11r3mnnX
ULF6gH8TE8/zu5GFXrE4BW++ujH2RtBh+8s02S0N+rHnseLpOjGyFoGgdutnN5xD1YQEaCbmrL8r
EXNQUB9yg19eh0Mh0LqTOnVZQWKLyPSKzE+e2PMbR4zNsiGllKqwNWDFlnwVL0cio0qkiP+e30sV
fnUaQtfcG7V+8zN70TEGMUx335DwvfwqMV4FsvaO3O2Vyr5CpD/vq/pRDq3hztXpHt730CFnPWVM
ix4eurtD+XA1GEaGynAulVBLwfoey+cEvi6B7FkPro+bHFQifLrAHx45Lqmnr0W3XbDTDxhFJcr0
ORSmTpk+w2UZkHDdj5V+MY8mJen1C0V2yNrPuzI/ww96XJzk2oouxFpUM958/s0deQ7SHfr0TewR
VrcNGnURzpnITo/Nlj9tBHhES1eAXNmKrmZlcOD8elsO9Lrx4HjYmUMlo6F0bUTyiPTfHzuSeLFc
GsiKtOARwA2MlYHJeHsS79+Fwl5bL9z2dMK85En8zo3JM8qQiln39562auD2nNG4Jaf1FWG785J1
XiQ6s1ifOOFzT5KeeEZ27bFd8BGebqkcjGtTNI8qumbhBGdFW+axMpn/3fwGdnZJVu2tKApaUQUI
YGEiv0u6X/LkjP3wCPJcznGfIChyEoCNXeZVcaUv0Q+FXcTWdGEOg+hnn4YdLHWPNbrl60VU/68t
pmqxqPSJU905s1/3pKZt7dkw3J8KkqnD/z8UlHp9JeaPHqxnMoYjjFZGUcQlc15Q/wG4QHPC0aKW
lnjuGkh5Xn/VY5z4B+OtcLmNSLPKKFv2kH6VuFPnsj1K5IiJMU2HWAK2vwbc3uJAHgMZ4jB1nr7Q
BJjgHthFRm7+bdL6sZzb2rHdAYFi4Dkc41eVwYUMhytOt622ohCqI0t4m+3nH13rhAYtYvsOziHC
BWwR7hdHq5WkECKQYfYxDxriJZ9aMA5rsQ+0FYmQxTf+BUMrR4iMfPvvKIIlZpbtvZV2z95mi2Q5
IxlTw9dF6iQtSCzEa5ucNwC46dwX5JOkJZYJ9PCvhjbV5snEYH/CUeuVSE+gs7QyTXZl7SBISYqn
6fPjluwvo2hVfHCvBj23ycC+jAqm/ZrI5wSZPaO7YQA3l66QygJkbnbA5mfnbh6vbrbZIBbUKHXA
vknbJlyJzK5gsqL4RbpXlh3mqXBbh0Wnq42e9HZ20D7BUf39bH2mS5Y5NFFoHEDB97RDPJ9+dHDm
rDhgJ6qE6im0dS2L/u6TVjCf2mo7rfUmEQpYP6QB/sBrdqICWvjK4x3nQlyeHmLmpZTOnM+AiAa8
1Vm5xEjuytfgVrCYEyyaCGj2miW33dJ39svzUbZqODj5oLoEeutJyw5PUtTIRYYZlgbO8JPhKxy0
GqEt3ELwOI393B9BD0Ur/4iA3L83/au7CyH+578cx6SuIqYTjP2m0598jEU+b+7/rPAwcHtGmAhm
KPsuMRXM7fJ8aclFVyvpC/nOJJs2kfbb+anMNEsOq14W5CuxZPalKj4azJYKz/rcQ70dfhWA9Nz2
/Yyl71PsSfxSPDmA4+wHGBL6+Nimkh6vB+42bqawbc/tpQ1ePOR62SSFROqUoTzcgYlezBravVkm
/+WpQiRWlWdKpmf3S8NfhY/Z3mH2H9Px2F30I3Jahcfn1ZYlfgBVFGYkserH4MYznwXLGxhFR7lO
vfx3wmcSwzUkBniC3bc4H/262+mo/EGJ0puVxCKfIvLfpdYs6zY23mkYABPOOd/Lr1j+aP1di0qD
RgFii4tiQlsLRMtduy50/Xhf5OY90X939jRsEJ5nsubl8SpAvL3/SXVPSkW1zz8b/X0wyqtYpUpe
URa4CFGm04UUs9IyX6FNe04FfzJiP2WERVgeVIhIxfhvHdG8gFA+FvU1PH38nh3DpMmav+nxLSGF
dQznhgSIiMj1roVtYEg7CF85XZXiBFDYayYjiSyEFY5A6ng5LQ1/UbEyrf6/taopLHGenu272hkP
cpFw2gNalOePObCjpfo0cJq7jnGsAAQTa7HNTR90+YdpsppwDm6+RuzM3LYasNwzjyUQKPjVwr3D
lYKS2nvae1yETXL+rfHkE13nrGTzRlKdlZlNfxy2GlLEGuZGMwJg8PfSMgXsA+zJDxQV0rOIkj3f
iCPg1Ok/RBU/ilYxgAhwyHBMV2/Swcmfm8Xf0Moe1Nihu2pcnCT2Q9jaaBAOHU6Pbr8biGTTgM6U
k0svAgSLRu9WhTbTm1pkE8wab/Do77qNjbpbyfSvnZI2DU+GMytDBZUrhR+nC605LUBIu0qa+NpM
sJFFf9weEsrhV5gbzgy/Y0s53aBqHX1EzCsxjLtZI4TCs7UcgiihxjSrRf6K+ZcxdkJuLIXZU8KQ
DHbCe6tnReVhy17c6BoLhxBD/VNErF57zgOiWG3HamkH/gMCxJ1RY2+/s9e29gjGWOecM6pZtcEq
lQo66MwGFq8JhQtEUtQZJeEAcJGMwWNpuZ+PKI1GbgU3OXVlQX6rFVkeYVF6c4HTUN7KKWFDhRo3
nN3fbi0y1+Mra0hP+aMbxIpysZd8/94UirsAdfTjogSDvKL98u9zktqI0m5oFfUbxk1ycjJlE5oF
Ar80lsHLTKJJSW/IW4Z34l3WWGPVGbRDePuLfwL4qWrOi+gyCX0pjf5xy+KzOLXhdoeEGjqqVu15
fENZqJo9YYJ9xsIQMwC5FdGhMQ187We8TRodJvU256n0nbGx0sR9/MR7LK8Mr839cA1oE/iWy/I+
FXfcLz8JpxA2IQkYiQKWHPSxJ2uTePAzDZbDV7bAhWVgDGbvnS78j9o+xcKcLblE+il9pTVyhvss
kHAyku73NRbu/vWvjpL35q/sv1C8N2t9voXbPAeYR3GRCARkFbaNamKZqVBndZ14z0ZqyimsNk5L
Sf9nbJxjsgZuOPZCNArMzuUF0cHZam65/OGQAUHaIsmgTbJxMFJ8VDHZ8bGQ2JsEXWhNTFH7hopS
5Oh/p7DU6STgXHohygczYwBwoORtqDIiK6IgBiLncbiWiLB0u/eiUeEQxKP95ezgPGRS5fTVnagi
0YEwU9/djj1AnrXaKvwQWKf/3rKPYK3CQ2OiGptYYujs4sDOjgMuQKFQEB1mBeZ7WQrx4Mr5Zx15
n5HBCMLJO1jcnp2ja10RtUUqIxGLp6MJiCntFt54JwkZy0ppz1e9z980mPHaHvifmPGcuqsnK4qs
PVyGEqBSklwmflMXesODcxD3VEoCo1N70nWQnbRi5AsnERJpq5jeSde4wj4t4Utx65IVQ4sHmDkZ
Pp5dAoeFuIy/28ZJXdEom5JWSZ/J+4GXfASktd9sBQyNMZrsRVgr9CyPuIbHftDYyoL4Tq949PfP
/bNCQXyHHvH/uQ7Ba9Bzbm8iCpNR24yKjRf7CzM/78dhuPCGYMfBqO4lG8fbCYvARMAbgdENGZ9f
oJqmd+TDySHvLjQZXhtzYIR071Ph0uAjc2LKeXllsquVM/uTP7s4vht9Wes604ByfWUAN2jeooa9
qtP1Yz+yE2TYWxN1uxEuJcMEsRohreOrdhz5e99A1OpzhDEtsiGOdZvJE/HJOiANF7cpZv7ipXbS
nekNV+OJHyYPbZs1L+twojUtbF2gOxQve/6CHhFMkP6ZYGV3XRNfcspOwzXRL6o5IYBwUAGcF/O1
zVBNDSg295Ft41NFoWf7gVm+hwTMvh/h497dl6vMEuVUz/xNhCESIe/6pTaolUzgJ9D2hWa6Ii5F
TEd2P/tiQUzO9Xal4jBeqO3FaKHx1tZHDPAr+55cFrWR4lk/H93NvDMpvFlrAEUVchg19ihv8vhX
ih3hsiK6LNUqYQH5M3Y+iREIoLRAOAeeV7kpwhHJRS+aW4rGsLyAHCCq27hA03NaEAoxWgaaEzgA
tCBHN4fQLwwmbKueOHhsAmEKcL/RqJKCrJ639BuoxTnXPpkF+SRtexpmsl4kDQlPnQTf1nCbqTki
zpSKRA93+6NMRVj4s3LikWU/k/LFJG6NWe+lNzMMSbcsdFpF/GgtyyRu2iEgVacTGW1RLn7v5BX/
4fNLKqeuqDoSHaJFG2di60AIsNANUSk3K+M/jxgNIPlUccvAzSBR49XBbxZ3mcmVFkoWCRcyov7w
WA+DQHyQs09XC41pcgd6y+gM0xhWBgXJUqeq4gk8M7mJ+82k4jT5hatBt4OHL/X4J+gUV8o+PTT+
wNUzV3afWtdIUUrO9f3yWCjTA/agFXu7PboF7pRV0MEK3BBz1F4ZxUHDLzKAlsg8cY+A34tT0I1h
zBzn28jKlIyhg6hzaDB6eCVP9So5oY76oNiXluabPCVSL+gDjNHhELl45gTirsrC8frqp3W/4gOq
x1kjY1awnNVJ+HrhiBRMZfpocMsu4ECUsU7D3Xfo+Nv7MUuWiN2MNmVcHiQtfmDSQfQaSv3Eippw
s/CPmq31FyUarcA7wKCnR692ih6xFjkzWrT2eBoYbD17pLmgSDJksvS5NQShWgmAbjwSEhsqh01j
DwHd40o2/sHGHCeIKUNIjXe3cQRgisOxDZlFeU6zqDt2HBUG8FH9LpXKy28au5EVhV6jU9Vd2Xcc
aXgEDCn6DhuxTW/kHRxykcYJ+JRHW768LsymJQN8xh+3J6HJu7FUYZWkJPUuapgTmIs57YodMQhC
x2zfx3rliYQfSz8laW3fwbPcBmv50LMMXm5uXJsCwqOYtGlxVMNqPBUWyEGVngFJpUK84IwTvSro
uWTD5IoNiLa5HRCBbYWb5gCnV8kLtm7joTL8zOPVmu6lN3IOjh+n0NZHWLNQMJ7E5Twz/Hipd9MG
XSFoNozEAADDTZzzLxoFTNzEwP34TFMQGhQHl19Y5aPEIqvIlAHGUTvfGjYDKmXPHxCPuuVxctyy
7DW7T+BRP3WQurj7d0zhJ3Rtu92CxnaMmzd5bCrr/X/3ryBFExxZcIJrFStoJbMuBvMObokBdwT9
XILQrALrI9/5zV8fH7EKfhl9koMKLR4yJezd5nY5LSBr1A/XRkxYhYWd2XXAhGNwcHy5VOO4/kPE
vO2KOgfZUGwK9njiS0PS+rPBjSyuzgQ0FTqaBdsmHWpoYbNnle8xa4sSpEhPTcYRVX/ch8VZVtIM
Ywm4gNWa9BUl39ZP8d3lToc/qBEDVRXiIViIpgNLpqIveE3/7ysBFuGzByeJCoks4P5TN2OGtHZ2
uWc+IQHk48TxPAMEN7qGV9/F22nXcu52pM8vR8VxPiUiU7cX7xgDUg6cz31tDXex6eOb8ToxsFWr
lUn6PHH9n3pTuH1NwTO7TK+Cgh57MPlzo+lkgQubhYopQG5xRyZFIlnTrWzCsw7fJL+uvqIUcM0f
zd2ZodM7iX40eLvOI5+iJ5BYBLatINkFoZW/9A0x78eLgiMbsNuX8bp426E/a4nAVDDZKM8os+yG
gjQJDGVCtBqWtePyKa9itLroStt2EllIR4sMhGSEiiUgGFaggjrP6tygyF0FQD0No/lJjFil8CKZ
6HcrxJabQeyRsvn7iMfVSaJWiEDy4Lce50C/lGaaYZ6ZntkgsMVlMSJyhhbxtV+XsqsWlslope8Z
QMEx7PSfqcLHXaj2Ogupo10qvVAUK1ao4POAH7peVazhMJNgxL55YMoPSgj8WUtGw/EUD1SO96FI
HRj/fhulS3wQn+9Ilutfm1IuyVFlbv2CZcFJPpRUvCahR37HpS6FrYY8LHF70DHsG6/jAECD26Lv
0e/hhQZd4vch9+l5k2t0j+jeWthRtkZe6Ygo0WNKSPh4zQrNs0D6B1sU/mISVyyXIroQiMHsTjMB
Q6sR+19r850fOMze6/INK0IncN5GgmPiGYqhjsD940KQqrEnCE8frBKpp1qDp/HmAlVLxZKtsXX/
VN/FTKW0o3mvoELz8KbEKcXbTXSGyAuOER0ROX3QqhaFPAOy247yvsEhIrSVqAUR+X2IvbqF/RGW
n2YlpezvWS0O6v/YbPQPaFNQUP624z/ec7nl/RYzXf58viWQWqUUOfmNc8BcPYHsJCJoTmLlH9IN
Z5HLKWLkDjE6DD8Zb5GMZVdsHpqarPB60ZdS4ufix5VyzASodmETNIpI77PV4Lw1Z3npVrdVN5+4
bxEcZvOQW6HBp+g0sYXOuGgmLcFnQwufjQ7EB1leXfr88a/Dd5+pyruw8LVNU/h0nsuALMctvUS3
U8qqJIbmggQ3xQiY1MFbFvixJ/6pAVB1kbr0iOHZ7I5KAdYGLEZuLBxJpngIo1lpY7EwcsULXWZy
7kDfoS9v5DdwUc6rzW95a4WXxjb4pATpo3BIQ/fazV5maezAOvYJ9HBUYlKzE1dVcpsTTpfppzT9
m5vCr7JOIj7kajATADTmp33MGmRDbTeMo4QSZOiKzRPCh+amNW3shTqRDTVtYWL6CllxxVl2Ua8L
LHoR0N7TGyHc1UUTzyZ0rSEAFnD5TOkeAAODYVcSGrifgAoBFB3PTm9zHghR2+hp9MQaFteHHjjN
yHBQYfxDit6iknDSj+EdHviEouWNhEzhV7dUcc/mdrpV3XUCSUExQtxc8ZQm0t2q43TB5NesQt+t
dlxJA52gON2pudWwDKvt8Ea6Hpl6yD5q4mm8nYXKAZuJ12Ez0peQf2EnZY9EXzu5keJGbGg0o/X5
dVbsfib/9MdKjJbYKxavNf5PTIl0t455st0jbUjXSHwEBmRMmpmn8cjAgrA2lQ0sS6cWh1HHToJ1
Y/LLBoFlsooFUICgXSHaRMBek5sKVJCWMSs3rJ8sxiHgmmNP+HPmOPr9edF/C82ISNka09U8/e56
QX75YDnPW418mlFkTPnAcPyYwYzrtDR5hxvi8x45d/3LaS/kkm2NCsBkEHUnsH/FXtDKYA6ybQvC
0Nvvm8Jyg+jsniznuXzUqa+daWrr+QRdveJwZf5HLqthj+5bno4K1wA0W2ygV04+iiJlGGrxCvNS
BOWXH1gHIYFPEg6dusi7jOraRYC4AvgrLavvEV+tmp5oaMgeGUeB8Awa+J5q4qzTsBLayctW+xze
MI5oac3an9oUExf2wBWTkkJ919INIyFrMKFAqTJ/FTse0Gd2hVvn20G4y2y0Jc6PaE+JHbFwwjao
27mqhlaHjHn/KWyDnULYvGv+Ntr/QeaCPYPmlI2L8cPhMdbbTNIon9PHhHN5PFk/S4lKhcASgHc8
I4El2TTQQiCc5sw+MwAgkeGq5VJvoleQ7pEX1BWwrx48LrO2zr9AqmIGg9mIjR7zgqsoYSmHNHoi
2m+DGRYgIJlCegO26m09j3Yh/gumBKAB//QLFPgKu2gOqtLbluawZu23r+Y6bnAn8QCU5LBzR0W6
gy19WXsKPsnajvzLEGyQYv6hgVgE/Mwc4D6m1g28EBfmSAfPyul+adhECODc/Q7Zgm8s8k0TZ9Ho
KfemwVtCwDpi3yjmtSqRYgiaLLtSEoVvp3m1n7rvk7LaFGGn6D0MRVhZZkNEQDdL0lV4K8yOP3Dz
NCjuabycST212Y4tEct9FKGicjDtJJfM71mnu9AEXNEqVm7smimHbc7Xh7dTXMS19Stxf1CvDR/l
XuwAUPPW5U7okib07i2TFmLqj2xgVZ2Y+p/Xe+Xib4Qe4aNGjw9m5KC2PDurkbMb3TK3tWqMojYl
elzdqZoh0XGXPHOzoOUfVphuq9GnK4Y6lTnCjCkV13D8BZKRH+7iN+cEug8kNH6aV6YLOjBTij7g
ybhJY9iC1XphwLXZUXkT0MGemdOexGwXd2GBJ5gqn5UbRe6XibCf35MAGBtel3ZAahIF2ZK+EZAo
kKjjFZObdYKV/TA7CmcEYx6GM00aM0UHOInLHeUJYgvoCIye32RNErAqICGrt0dOAXcAjJ5nmvIl
02/X9BWgsInW0GbzLT3wLns0G/ErMohZGv9Pcl5htRMadEZetuL1Hi2wUQn5MNWB7+0dTreypQ9H
P2ao2md3ILEuP1fvmaBpK2sjsQ+tNvMrGnYPopu356Bv9MEmRKAsip6d0uzAtkfvMr4tihUcx/P7
My5kSvaOLop4pjtpRV37BYfHP/VvrGk4OSjKScqiR+cR6J8sL3mLAvjFDzyTgLoM2NvqH3i55y5H
P6HOTfpVrAlch2skJuGGsSUHf1AP35+BA9aerYF9qvza6lQMtByP1sTABYmDw9ucgNRSYAOhiWvO
P2PWrSuZyE5SNaLiL0JtGdUNjSdn77lYw3FozjSDW097PCvBofFWAL4hJMUfq8zCC9f9/RqvDtr7
5LhlbVH3S/cZiHzEPB1fTgjf5oJnLETo/+e9nO4DMTI9eg/Fnet6rA1to+3OhPR1NWd5865QjVOr
FVwogn6AcARlS/vSNbZljtFRHc79qJcOijbqBdbfYtXXDaFyvzbAHcEA/1ebjrlq9BYs3IOPgfEV
bPMgc+3KOWq2mi8dTe3VIwXeZCMUAmzFi30DzK63nwBoMcKARapjNub8YlVCVOJ4HqQxeZNNdJAn
OePEu2tkZAF3JdFEpIqOCE9xqbqEo6L8wNvKrv+/9vtIt+tIKvFlmJqVO32oSkNQFUwWoWYQXauw
Yqhzt70ViaaHUOGtVVXaEBMcWQSm5GN+vToVNjiEUr0UBBht+ldgauWEW+ecKB896Gdv3pMIcL/6
q0lJobSTPiek9u+QSmSGiPJh71RXEeHgfJH4PwiM5MijYqSC+KR373qLTyUFzE0iTxXgKcZcdGAq
vu1hB2+bPHimHKvUISfneWJoqtie/Pom7n7ysuAB4eF6YCTwnGzT/+Fspgj+a7zlHM/V6Xu6UbgY
bHwBLBXg4n5LuioOn3CZDi78iaIfFswmEMwj/bON0zMqw17TMXe1Tq92IJpsJUInnVLUHcjqWQ1g
gLpvPgwfugehJbhQZ3iDLsteiflf1BNze2RaFUI+LsK0hVd7T5/HL4PYtsH/ExMU+PsrwKj6C85v
4ihJWETe0xXf5nCt/w6S7HP5iCg//23lr7jxrJMBCBOeM7vMEKiihSbrHIML/81WxFs3qkzEh7V1
E4g8NT+HzZ83TZGyhjeiK1anRh74OTY9PwPSPNIIAKFyX3LCBRPXQMDsXa6DeV+44hDiDlCn621e
UZERPJF5b/M+jZVsjZ7Aa9PPfVh51nILGQiy6HyNchKDRH6BiUYIZj/VpAUeTB4PVXYtLH4jMmx2
VzMsGkdyum8OrbG8e0vtOMMT00NFXz45I4eB66Uq7R81Yp3FVgGit0DCZ/YBjL/gkuwlLiMCc9NR
4ZDviIbRo5gfYnwXrK/PnUIeiwgbkmGxkJQQ956KDoQDrvPoHtKyO3nECJXFQYmFaN+QnACBVpuA
H8obZc98gcGHv4Iw3CC4jlVBpLNAZYYwxlir5tg3+rUrilwfedJ8F46bPqDwIuC9MclLpzjGH5ct
kNCb7MoLgz9jgxtXXEohcJySwZe8LyQ3iuhHUXNe66LnJLh8oL3GXfuAZw0E7K4X6TvxOK3ql5/8
O5oMUxVlmMZ+MusLM09wQOMEzJJTJeiXheomL/YVqs7v0+dkkAcAyZf8KfQFYmFaaNKffXt4ZV9M
CWlESrUjQ0ekBPsb6i2wtmGNLa8Np0CL4eTPVXCggJ5pkN7eepzcevsrK2L4iihxAObdV/4js16/
IFokwL5zoJcWUyLd/I/UiIn2VAarzrjRVToZzJ9ReLD40iEDMyuO23SNScIgEpCRjTJe5szz0ocP
J0iTx9yOSK1k8tci+MAWjT1e9npBlxmeWsiUHF4qjKuAVZlmkI1fu83EzRcVg2TN4AfZCUph86PP
4FEP3jVJonkqsTPlpl9nOLmKi0qFmt61dNKmdUgPv8YYpIHd2KjUL0pt0y4sLUbSgCkcILdswP7i
aMIeXN1S8PffE1F208B8BjXtybYqX6ipQ3BNeMeqC4dgIdNtdU9b7nuD3CCYxEekKsmuMB+5oozB
NWhk8S88xS84e+RYUp+L3cQgXJbmAgw+0tMx/pI4n6wnIhZ47RhSMxqF3wckTwiTQEMwfgiA6G53
OBAcpZTevsPFaW6PaOgvhgfwmzBMwvsXimIsQG0cL+LH9KOLurOuAi8eTSZ5/efurv/EX8TQLyDM
ZF3ecirdwNrO0QfOi/aeQP3PpcMk+uSfBDJPEvZ14nqCOSgfO6XPR3ekB4ylKvT/HHp/YXQq9pSJ
QtyeKbRgfRpc58n3tXUI8E2H5jPp2U2VOv6nSIMVqOYKew3MpDREenB+9yDGLcrqjdte7MXR4Joa
J1/iGyZeZBmDYjPyq2GOFMTFgT06NvQ05qX5jMgiza2ok7pA9GR3MjSGKCgbdvog3ywP7d38DP7Z
8C6KNKnoL4aB6eoPTBziBziuD/e14ntX6Q+io8oILbXdrI9n7KBfncaaFILwDzxZWBSVcDaPFJ06
2R6MCMI956wpItm1LPZSmfQo1T5ohCNDEi/td1PxMXs8firRaOcRkYCGp3MvSPRHTzfZI6Iq3+Z4
pCwDP9hCtnGEFRwKDCcgo1RQNF5UMwoxAIYoGKMSVvmMv+ZULvt+Q4MFfkjyUQ4fd90ivwJh0DBE
0lFLIVqEk16ADxFU8adCQBhBkaIK0yS1TM7e8Doh2RsJL2BY0EUO8VcMCVl4o7yYDHoVfbGJBTsn
N03wb50KQsrW8g3TNbaAG3sZZOmC8evbaWUJaegBDZ8x1X9VHgQLysKvYOhpTh1CspqnKxqFalIZ
rPnmTl3NNk5nbbo95IIB07UfbeUnaA03rFsc5pi9qMelZa+W3LFeg3uRZpLQw9ZyUwJogyS6hX6h
TItNiL5+KyxYf3BDC4y7zEiblX7XXMx8Yv9dyyHG9rACvjc38Cx5vzFMR2IqZuIq/Zgg/cz+HB41
MtJmaaB+DmIyvg6TvsK+i8926NHguvc5D6wUdNcV3r9GW+6AD6JNZ4adu38Nr5uSbU5ercWHUx5G
4gVX4FhQt/AsNn8AcT0iGRenNNKyl/5gNJZOjbGkFHjNNS1ptSiKbserz1MEvQwT//0ygda29SrM
zoHaApAgwUt3KQhby2/fCbXolxnMghxNxXjGbaJW/mpG6zeAQrmh/bMyNv/QsIzoAV+pUqq8GAkr
btx1Xc3INdBL6NXbQb/2sDMCpUWoOD6l3tHs7FHL9FuH8vXAb1q65e4QyPcMiWMun0615Rz5Cuo1
LDQDOOVbgdFg6h/bCaSefavpQf2pMQv5k5BAMorruSVX0U/dCPB2GNB8K2lkqcdt0tdwxyy/3syE
uh27XzfAxQJxn2Gra0Z77ux0+c9P6JZWPoImPhvPUL+hlG9rkJWyLtEwVQzSJIFO9gk9Nd5x2aTU
JRWI4nJJc/CZqdKlvxh33qlgfKSDUZZyRlQKesGZdDIrEIFdyYsw1MAouq2AkVGK8yuZQ8Rk5chM
tKxxJkR6PuOBFQbRl78yEohvCWIuypGVM743HBHbFFgK7pW2Kw9/HYGmxodrqr92LEzCJ7DPg6OM
zI7HrvIIn53vABQeRa91u1YNojq9dizph4H6TlKh9Ur1CVsS6tKoyB69yzln3nad9DU57PxnaFxM
vLuz+9AgbA4PvvciqGjmi0rit4USBdlDKDMWsXhtFVWZMC0wZzGUOIhcJwbNxJ9QoZMKCTJKGhIO
XRzbyq9EdsIoOZOYI5TuTdPzTjY4s+CRHWc+Wp873k4TAyfXzZcHKqRArFje0+W7hIQvAvqlTckV
hjbHJ78P5B0PTECZ+fJCrylcSHOmsRW9lzfW954QCcpsD9Y7QkYUseH3vgNdgIpIKv6u8Ez0fqB6
5etDtZ9w/nnL++OaZFrbBoDg4jHOQId1Td51N+slEU3IWL65EGQCJXgxGHo6n3SpRVxAYiQYx8bW
d+iXQFWwDK3AybmbIx01Hf4ng09PaIZiJttq95AM8kwLM0nbx1CXa610kvV6uXe0GhS6HoBflOQ0
EgQb8blLBP7N2kWGjthd/6REyxZToalphDtsAEb6P5A7JLZ6ETOp9sOtvv3HRphB39fRe3tKkY+f
2/9SefEZBYiqHgPKpF4rAfOyyjQEZpmc2IbWbVfju2l9Cu3OKK1V/5zkMePRANeTjYy6T/4Rni05
mHztL7xCeIDP3rmvaQz3Zkaoldfm+RHlb9BXSJHhp7zyQQKRaFIRHnHgrCbMh5KHge9EUeLbnrcp
VMS2ok8BdKxRj6P4nblam4kL4zdgd/rGD1L28ct1yzaXWgaoRXKu6XZn4ScY2myJBPqFgSsTRCk1
gEeryrp31W3hqK3YJw62rs6vv+EE8pEcMuGwNfaDjXtEw6tHg8Qs+60cP+FJfmQVVTJuzJmc0Sxn
E73sXl9vyUN/6RSUZCZJ2KdV9i4sKQLAFRDrWQRAxKeJxY7EPRwv69nq4zQysjWhLGRFEa77LCb6
rJLUMk4xbZXsamKixF8ya0MDtL+qRANFrcili408j9/kPEakh7VdJbFXTtUkypGmWZ4Ku+y0AN2L
QT7GiaqNi/nVSiX+Ua7TgZu8C1cLI3b21RSw8uJ8vTB16kpH2JvKTTfz+ogHOusD53oIsT/srA0l
mUwnFRC4iQ1dA8IA/oGtG9ji29bBndqXSkypGfxlGUksM60d1eU0nIWiu6/ktcuka4mkxdwSW8L6
Bs9xaaKtoVtOnqhvI4tFekSWhQTHnyfD97hmpk71IJyXGMl1UHlaRzJR8I+3ydi2pgha3alNS2a+
cWKhYy/JcvhTWy7XMHE2t9hadEf9L4TplOv+ANHbDgJYpQkZnDFgyPDK8zGA6D0rwxpa13sTmBh6
jczjGVw5XMln34fFSAvNTuraC+F5KL1d7qQ+IcrjYQPjfW7atNi6IKIBRN738fc3oy3AB4+vWBfU
wjRXpsR0NloR4qpwkSjDLIYfyWdYZnmyMMtqYCAwnsgvOOJIPmPHBMMjyLzQulAxsM/BZ5zN64wY
QZFhmHDh1OEBL5gCuEfTAwEqQmFsHDIDSgMepTlavw2rzlyrqnDmnHyYHzIjq5aC3NZXIdcxeTkS
PDSWUB33O89KTq80OZKtwfdAewL0SxjWetu/6bN0NpzW2xgNJKanxx/t9fdRFAL89gBZiyz4955X
mImqhZqdg+cyAGLZM/TkEcW4eMsIY6G98FqJO3Q/ad2YFFEzUo5BlJYxg+WJgnkVD1XH4cveTfcd
fEyW8UCHXkikBfQw+6yGzrBvu44PT61XsVnK8QEebS25PEnz1qwSRMwXjxL0LBT3UPbDuwufzjJJ
hiqXGSHeQvkF72ZaRI6t+brPiyFh6pR3J88IQgI1+7U7PWcqx8+75NjSPNEW3BG3kikr4U8226kP
iq3gxTvGk6B8Ii0zK2vI9M0H/4pn4sW2Wr4o6ZN+c+9RfeoZJhQB5Sdiq8K+DLDC2bGndQJ1MW5m
8thI7NNvKWhKK6kBu0HWJzAol8RlmwW2lrmRt+RUOmfuY1rI2andhwOAhNvt8SN8AR1HJfo9rTyK
szlINN0ZyeuWGoE5kAMzVPGBGF9l4n300TRrf8swloVGEkAsCxjrAZOnSGaiKHsHXscpPxdgzFRI
vtBSG9mDnyEXlFMTWER7ZI/yagm7xsh6igz6DnS6ggkh6JqxMSYEjRgr7DICJcFpv3ivHsXlzdaY
6+7Uk1HtLN6hxkXxGtaEzp3St3C/VtxjUs7FW1QSs1GNFha64wGdsjJtVCFesYZ3uZCWXo3Dq48Y
wozK0/OoCA9TxPNPhXOU5pEQFKLtG5lzQxCcjd5iV7KQEnXR2kszUJfRweS29AMbWHLlAw4KCjqa
v6nOhfYFjtiCEA4c/XSs4Dw3ql/8QdLbgcN0nbAAqJej8NneKWa0YfDUTbaNLEEjBmpPskbINdnc
HeQrucbQH9yBlVBZCackj6aAPRsQF8nZrrtGN4N6A7WvkP2PtyWRQylu3MGL48aVzrt1Xa32k6bB
F/0NCMbyWUqgdu+VY/yb+gwqLkNPr2ujilcgEJINPUOBwhF8LBJ8eVJRE090uhjOr20dP235pf2H
+y1qWB289UZ5nN3hO8w3wWRbTv92V9f5ByM35l5jpjKqyJq2F4sC6KS0/izwGKdsLg4if4MG9ZzI
C1nJgRjQZ6a2Dvk4CdcDM/Rp7bbM0dzN0sVNvGx9n+P1KbU+huMvY+PSQd6h1XvKgwZazYyykcHd
bT0SHzaQRttYDqFHavE5+oMEzuZsv/pAZgg6i2Mnyngb8nxLNJnW4dQBhTkefdhDzxM//28oLipp
otlf30iKbzGgFlHxSjdQaVnXS3nUJv17cDh7UNsBenF+OR0RCVAlvbIAfLux4TzeTzRHuR1JnDVk
0XXHUJ6kmhCgox4XsDowf/eoZJkvDkgmTsPdr6LBU2e1DcNg+bnyjQmqPW+CCivztxCN20MMskG6
TQBmDzczATnhOn/4z2aFg5jlHFErEUkaSIid5xIrZ/xo5vflWQjyuoiJq3PbGj7w4LxjzCvMHZqS
6lAcy0Q7QWVWPn90jqqxbRvHGALwsStfFogPSmjEQpPHBSQJ1N88UhakdPuo1seCzo9DO1GYep71
Cz1Cma0+1mPlHNxtoAS/Sxm96h+Z8MgctpbufO9im9x5ECOEAy6GRqQTiX/FGCxXVFA1O5kc5oeg
M7FGwQ8KYWbpD75I8o9hzWB6ikrLMmohwoVzIESP43JfIz3Pbqrw58gtcv71FsAw5jTSyg7r+Bdx
MXfMiuzIFz3/uacUcsX3ZB0oZCjunN1IJ1LJQ3sEVSw1qdXdm69hJWOd6wCxSygKs+XjqgKvxzGc
9F10X41lBdV3RW1LbQUsS+yXAl8wDYj8/5VH6sONRSUrX8JVhJxZIRC0GV/QsodV5/hvDXL3VP3t
nOrTj5gkKSNfLo7StyRnLmF/IVSORqqsjnRY0E9+E/6YY2Quf4BZH2IkoQDXW86oZJCqyaE1ujA2
LKJsXw/ORSb0+ADrViVAzVQcHaJjRcywNgqVLsG7NqD6RR0jc4o9FSt8c4CVroLnzcOcJ2Kd2pZW
QI/NB0ZA9WSOtdQDuIHkCCmm3Phtvg9wvk/U48Oh1QWE4i9T8an8hlpYvUwRYZxU0GLWMKKYxNYh
PSs0yIw35YjdFZzE3aGW+Mb5nBdM4cnH+H2XQTbNSY2GEzMiz8ohsXVjsF64g1SfcPeJaKLpR8rp
cExS4Tcf65H3O1aAOFsfirzVxdVymmUsAwDvBBvZD2249QHJAGlc7y3IxgJCSZpsl4Nfa1Xk3kUH
vjFKXHOtYKGrjhnMx2dXAhJ2wFK3mGpaBxZzRupslRQOTj613oyVvH6qi3sH/kTv3l6IS6DMhxT2
M20QAmNio8iRwYC84oZ8uoyXAXvuMM6nYNboCqP/zrEE4xh8HSZTaSDV97zxn06RGsAEoqCPBwTW
8DosbW/l9/aQOofxFRgio5lbFHOYgXZnwKnqlPWDy7LbCa+GTjPV+d0QIEqP7m2q9pEwaKwfL+us
B3y8T5YcBXQSBKy5pyT9ccZbpV83SVD72I2M/1qJn2D8lWAj8aCKbgsq3WUlOwr1lubHxnRxS/3/
55tZvsdN7oauCxOimL8ad2WqaisP5/H89w+9rxrjvPQU7Op8iLKmT7HqBGcf2CiMPOZgnHzOG3KI
BG9X2rbYO/odDBlk94IaojE4LHS7IBKhCHSAlZUZuYs2Zp4+qwJa37qimCn6/GILYt2Do5kqjW0E
VnMiGJi6a7JA5duN7MWdWIe+v6PlqWlo5tuUgLiRb9HBYzIQwVsDZwvukg/dwbDAh7xkxAfvY2go
rL9zh6dHDmtdUMl9AxnKrjywzGTCR8efQA3kq+4M0f0F68kETxqm6UjjMCH1Pcz7VwIZMrnw0B0K
AjjlISRCXEWvURegEOX1Caubt3vZ/6LrA81qWGRk0STrWBs8sZ8TVpl/8Bw/sPVgxcElkjOPerWk
wQKZIGfpGbEP/3ps8sobco1xJrYfB6jPPkw3IMXwvWbGkcEiMPwMCqli5aeFOuixM3obzdf9CSTB
3rtnXTEdTbcZpkTpqJvYuTNFqMbqdZOWPQJ/MwB3yMyzk6wd3EWS/5rIHeaie6AlIYuEOeWDGJFU
ijIdYfyj5XnmrCdjELD490KUb3tGaU9OnIfpzwostHlk/zy4Z+UAopKNuPNg0XsVikMHvT8fqgsR
MEwRUATpsuuIXf2nX0Afi0UKhTA2X87T8C64nnWB/RA4qeXH4m0lWWmvPIe9iDH17nX9yiUBP/t+
LPXpuQZ/W3Nm0nNrj1x8a+tJTjCCH0sDIWpVQg/sHNmCDVXDr0istwKfxSIX6yeid2BtaQuVncuo
r8AsudagP7mGlUQIBdAsicvtVJ7NtWsWTa+iTPyZ+EadNoYTga+vRD7KKPL7rH6xmY+7w/gbwWFQ
7kPUyczA17doblWFfloAJwb1+LM7civr3DhyC8hWEXDqwepwYBLmZL83Hk280O/qsE+KpGVChz1K
5EpRWGrsUH2mTDeOhGpTP5rEJcgMhPovtqgt2tO9559ugRnPVdpB1UFHj+peAkZ/+Z9+yBN4mkyy
Q0Zm/Snzj/TeCNtR4ARoK3KBuabNti3y2bOkH+Nkcc/9FSZywPNgTNz7RxcqfkGYuKMvJy9Mm4II
imuAQIkFuPFyaW9au+xI3cifG9l23GzhpWcBCkgTeaZ55uiuyWLyVTlUqNql3JQwOsDokclEXR9Y
JlzUEPU+EVGepO6IA7axloHP+IiHhrwMJI+whrE2PTB5r002PtXU9ir+kIRf5Gj1xOyQDb9ZQUm5
wu8TPTSeA7y3Hedob83dkMLkkaO1G15mUFMxkM6pdElGbd9nUSUBazGOUgH87YIwM9KidsWP17C1
s2KM5fTdcNzcKTAMFBWa3O9qLKFZegkbuY2+ppnZfkCsjVPA+q2nTg0sDCi+cq3SgFl7nUrrK+0a
mszOoIrRlMA5svpqjXz7zX8e4hiAUik6mBGEWIenDxVRnnZq7h2arjpGOJj4K15kZVoXJ/DZikb6
eLCRFQoNedc3CvplTdjSSmjNZhCPOx3PUdsj96g7IS6zHNh9Lo8qRp+sHdZXX2y/bpn0A9NsrBLn
LNnx7hqf5EYLj3SaBCBJDHQzOPWtEyBnSdFLC177Y6pJjtkapJWlAhUPcPC5D9ecwzyo95J0uSYl
PgMrTmlAiZWr0FWylUjQN4lbVHI6QEg8+zT842HG2dsRdxIcgppwJ7fi6hc2ZUTVLiI67xDsUAx8
UQXp1uAG3TizI8AlCBlXRJzWx2tXsGAl0aLLYp/SVoIM2d4VUWo6x97exMketlzjmSZdBbU/ntGC
T2a3C3Kpo7ni32jUVqQgd8j9hx94gukzuomy4+eTQpn2WOVvaCO/dLN0noCpE6s5ig7s9ETXs67Y
EAHlGBRZGyCP8hanCS/dAhsEebguzlGTOvCXTUD1vO1zIM0hXzoBMGJG9N+W4TyxAUzQDllbvSgN
5a1keM+9Zs2pMIwgNL2yw2FIdeUOIRPexFYIe2BA8eRFgxTXillVoYMm09FSPBhHexUSSLIqAc5W
SXRSLaIaVJtbuF1c/mThdDzdppvIGt9jcjGm7jz9NYEbT5hzBkfR7S8aOJylj/+R+ITfzGRmC5V5
Tq+B6hg5AGrCW0Co/gNSfGW89Eh4Ag/R1HMmQf6LcMG+G5tYhigabvOmilaCrrIPKtWbkFJ2f3oi
p2/9xOufapMd+SiyqvXzRxr+WKe9BMxJ+QaNO/d0Zczq17D3SlZx/R9T47NJCBjzQsolR3Z+ZheF
PbaeFrkntsJ6bjFvKKh7lpjb5SHOzf+U3fNB7pCABjkj6/0FYgNKOzlQ1yRNuF4GHdx/zSb1mDwQ
27RWGCXZ3b1SV7nA8OP4VTTgD0OS3+Zx93FmOgNfJg17mvouhiGZwSxVNO9/QWj4y6/KHlfPHU5f
TVujTpRm1xhNNVnsj8G6bJowMkPZz3T8qtVkSuGz/w5mCy7sTcpwBniKClHXLyCUG/3rHwVj28qH
K7J8kRt9YPTepsl3VXq2AVK8wpGPeIgnPVxmtvMq8IPT5AnX602hWZAGukC/NgsRLQb9QBPiJRM6
Vt7WOKkA7lENuOAZm5wqwJpumXBbSg+mxdwb88MC4bOXwSID5eObpaZVh3VpGCvjsVAxZUno5aTv
cmHM6R93jFQPXttmMaUifQrHYOe0u08IU55RM2+r7wh2r5w/iQf6sAphTXiu9gkll0Mmev1uYTbO
W8ze/EmFBX7loYFRgiAiJ4OJgWMfT1kSG8mwBCZMR0Gp2VXKrLmA2ZhxrhJH3NUYEGfYHGpNwwNt
COwThkv5e0tbYbuPBV0nKWYANAaorzgy2qJBMCzVrIYJvKrEFbudW9CrPnLRTiS3DpkALtFMd27e
9QX8oUIdLDQCI7jCpeJJDOePXkDQ5G9OS5/BfC2Ir2RaG3aJTFncZP4PL4bXVxv3wXBjBNzD/ECy
hPCn5HORbLaypAsGWkFARrhLog3E2D/yOhdCthFCH/PfmkJNB40pVvYer5UW5bcsINd3OGqApi30
1uJxzh62/MZashP1Lv41i5Z1AXuK3kuCU3u1Id9yVU4r4nLik6uyoA9f+mAYmuB5h99c2gsjALTT
Gml+l306UlFBj3LnI8W4p0ctC8+nz5YU0f20goBS7S78fr9fRgN4Hyso8CJ4wOpBf0fTi+qnzkzY
pm8OmEul6s/tbGkci15hcH1sG3hMxvVetEtwv+WNYhkN9vAhAdqjz6PYI5mT4WJ/qdZRmIpVh0Yo
lPJ4u0MnjCbuNB6lun0JGIk/L3elmL+imOngRhE+LQNzHN7aNwRYOKDs+izlmosyDQ305QBeIqHJ
QJgR8vHsvf0CnH89Hzzd0dQa+tlHwNHgMxd6wFhneiH9yB1z65KH8gE1xSLH9OPA40YIqnsexvMz
NkOXOXdV+Q4AQ9KY4GCKEZZ+BVfqef37iLCg0SjAJmsz6JJSi3UQGlgZ8WgJSWpZmTQNExX3RKId
n0trOpSg2P2kQi5eajVuLHK2WHEGphdNPP0AnzpzRa+ctANZrtpzW7g+s93tuIlTZeEIVTV73Ej9
WWby1HxogmKs9aY60dFB4r/Vg/4dXUoGLcW1rVT6I6llHT7zr9GB9BnQ7iDp1PTpRYb0B/ged49d
+rxQrS/lMcRSd1ezJoBw5hHiHxpB3/6c7c7/bFoZ72JnQIIgDnuxXaUNECzevJ4lqOVwK1qgDXPR
tBg5Jq+EwvAvXCrBBmWnrxTAHgMwtZzF0iz1SFpE2voa8hne8CW43VDUO6NWRTClFJZlgHlAiDwz
q8oRFnM6sHJdmsQZFcqZomMWbOyjTQv8aRgTQeY+ycH7PudWwT342mIIMkqzcsMwEZKHkPvuk+4A
UQJqAEQcakFhkHhqLD0VtimjAWL3r60w/Ea1oyp/bQaUWjrqrGpRRX07JSVdHi/GmarcyQXQhkcy
KnSuc2CdecG6n8F4LRJlSLH+vtPbGBbeBWZaL9IF5BHgsEmKKamqQRfCIZTtz5ZuZACXYLB+KSks
DLtI9uXwnlZv5Sg/2sZ1yTbQvEAft9Rjq/QbNbrbcTsh1MbtIGQPDhFJppGME4VDohWzzpVWv3VY
keWoyS+Ayq/AbbRVX7UcEfHMmsO7Ba4Xxn/RgIjt41Ugnh+6nUZGY1l7TyTEpn0fZWIcH+5nHQvF
IYDLo1psfBBFEPIRHqCKax3OdqzikqzSUrHNHKzJyhSfVXf1ghem9Lrt7Hv0Zht3aba8d2qk8Z91
jx5tB1mKyX1so8Q2aZmaYvxmsdGeoXbz7UNSJG8QsItljuaxpiKx2d4y7OwwVnlwoE4JnuI/qmPY
EJ15m6VR51Q9bFBV/LOXrvYNBRv82QHqKl4/WZHJZBN993+aZ73mLeFJUvI27vGW5KhlamW9Mft3
BwW0mJP4Q2mjqaCuC8p+GrIP9LbsIQ8i21c4LDW0CKA98tu05X4TcLL/nDS67kgj1YMveqTh7FHc
TSpVKGAdk01Zm9iqbSDoO1lBXyEvbldR+8yqi2R0tG9DBo63AxPX9peG92pUNdJjKNF+dQzqf+it
5d3JkOv4+BXRTKraOE4evBOQQVmSJlWHtkyr21esqbuDml3GKGebwZf5iTXSvV+57rv1TLz1SD6c
EGgi1c2s2aBMEVgTOmc8QTEVDywVnkRaEcsU6wkpLCvYrX3qp37qPyD0lkET7KSRVfJqtHLAadAU
uGFTNTuqPUN97XIacTmuvX8Blq93PuKwaforhydgsN07dyf9My8GgJrtgwIrLnhUldcAyFEDALh4
30JheDf/MIj8KxYL5Ujkr63Ks6l+wm8YnBRactDRVvMH2VJ5VJflNwX/oFU7900t06zMz2QJkUwT
Pp63FzT1a1FG5RaeCvyP5EbtL6vUDKDNE5e9FbnuM+fTbvemzfgx6BC09hxWX7lEJHLfidM2P90N
s/xenIh1L4oBTmClvpx3Dgkb3TChXdv1RP+ajXlPvPuzBf+P4IX0QOxClKEoYQp09Cy491E5QWmO
da1rJ+H+T8eAWpKt8PaUhbXJ/Uled0ynDOmiB/DTvIM6Jfj1mIASkV2UEm1jn4qbZexpBq+J+Hkr
jVjQHg7FynUPdjT0btfgv+CvLEhXKioH+0Ddix7G3ezA3rvuJYjhqlB/7wgH8itFJ7rprJduuDG5
95lMPQuN88SiLcbJvpSEa0ekqenLcnxhDWcfgt+hPZcsOlMv3jhsVVkGBNfEteeVNAakZxBgXs0q
srxpyX4fzP2zaa0MUMaOetdVhjkDrJelH87D2SDEFlwkjn0nhnVOcsgtNvDsbzoBxvs5oYzCFfaB
2l3fOICJ/v51q6sDS3zn4stq4QRjn3QagBsIxw+kKwQpjjKhiOfPs+wqIKcdLto3gAbtHfr6jZEf
MbSNQ5yxFQuF2ftMz7EIDT/lmOURlLvNJhLmgtYDPXDplQmIWUFkpm2JE6ubD5rq/fOSTN09r4jU
rLd1uKITFyUqnpV8Tl3PnX35H4+gMsEP9eWhZ/APpEu5GRpBkKfgjazEZtIDHlFpMN3ll4efz3kT
MGIGp0kkpVuO5WLJXaBdEKoyxNc6WnR+8Op/spKDWA4HXgNbelnixHTj9QvsW1Lnf3cRQeEwbq3U
fCrd1N+9uK12l6yn7VTY3MdV4B7oJ8YLcbtawWG42wXAevyLNrvCaN3qZakelZ4d5jIOsBmWLLkV
oR4/egWcIB7moW1MZljEdl6dE/BdMRouik0V+Nz34uSpASniPryjKixhr6OcGD5UD3gzKv4stYFk
vAY6Br7zsODJs6KsfLH3sm9EK7vjBLqFxm3WzsjDHCVSPpBYsbMT9u79HNZ6fTFxOC4dR5jRPRFK
64Dy9ya8KTMEOly/xiLnXRUtSQkGAas4gRY5zFEKwZhk7yknn7irmYZBrZ7c6elRWK7/ERAu4aWH
9lDAJ3leTElqeGue9jkEmLwJL/kOdHichAKfInhAGHBZFJ67AtGCTBUfQ2S1ux5mjNWmu3Khn9Qt
hXGHXczYnuwBF7WOshyYnL2VF1mb/wKlqfGEhY8Xt22elPbWqMW2xdb/KyHsSAn/dkhn9ji4WfOX
KZ86uhe3ZGZLs5cNTtZ7PLsq+zr83ELUqKZKnSCaejY3P/rV45fBy7tyUiRuZd2iCavInNaE1IS4
f1LHC7UHLxPPD5oyGE1eKC3zpILoVI103AlYiaSJDV8I9uZ6SBpSWMIK2UAH/PBwCu9cbTgvb/CI
khZsM2y7ZS/8skl2NuB0RTqpsNavwANEYwpUWy6G/EUnc0/MwYpVEP2wHWX6Hsscc8y/OGNVzrcE
PlVKz+fMGyzijUYe7WBCpdFzGn/7nn9zRYLF4n3vHJWjPzsXez8CnUGbGOk2z5FKAWrTenlOzihJ
j95C8aGPuPXfdW3E7bx/ras3XbZVnwVNZBwT+NymV5VFTD94HP2e/GGRNxAR87TBJOAwlpAikkQq
Cg8INwLA9y80WWtzPO7CS9oiDA3Q4GnC34tVa0FL74tUfTTcHvMLc/UrWvJnH8R1ABBrjJk7EjgM
yfGtQIlANwnHPra64/cI+LFY6UpSFP6qqTEdAV44ihbCv6Bu1RCLLKpgcPDuVhKVRks/W7VelDff
R30esoEKDmct6qD4bKSN1SIkUmkKX3vigHFTO9kJOyHUBWd8kO/2nGvPFK4P3iR+Zr4N9MAZbR/p
Vn8+8YokbffWF168+b1OAMvmewVhd3F4qqEKvU54/xCP8VEJoUSi690uRjfIFHRIizcM0gc/Ube4
MhpMoEbSPsdsMDYdoc177ndZsgBd5vz3GNAvmLIlDzQqVhJKf5Z9+CG8DMnIDK5yMLlBxbxrHSf7
LvXbum72YHenehL+y5plS9vDke2sVCDXoqcdCq/Nhg/C+VibW3B8nOafWbbHFfU5BwKXylwbOisX
YKIMZJ3eozZuHTZ7KD8PDItS1k/NVJgtwmMyVnO0TphReOWzE9NNJez+PkuNyn598awxjArDbWsb
piRlgri+vnb2M565qsjsGlBP+kwb7DTkwBfsFO14e4sRflnptlC/XZyZwIlBGogLd1mQR1B018eX
s970X7ktXbWggnf8+O/6lZxoDWG66R1rO/h/EXiTzar2zJBIPy+qbeljNV65DChjjFWhD2+N/6fi
5XjxqjcaDrukysvN51cLrbZPCqmkL9Glf7Q8TH5FPaZzgrOTmElRFkeFec6d2EUgwpjh9S8yCaTu
geifiLzMFu4Z0o1FZpnLZlXIqz3+xNR7qmC2QAPit09dW+QFSQ/8/OpKctr24d1soo7V4RXLljZq
tTjrtg43gJiKCULrQK3FgUItF6+N7DkLWyfCfAoZOia3K7OT7jMJfB99Wmivm5apjZ3p5UWAkjyp
GNU87tkcOW29fliQf/EGsc03HBUunqPE/BsHxun2KTkVmy/k9tMrN3uUg104RKajNa8bxSuRh5Do
cMA6n5PX0Uyykd/i9Ut0ApcEe2VqMRgBDuaRX6l0ZaeMq1IaYe7x4lG6L2jrijPp+x2ArfN6qxG6
XfVE7e//4kLMaPRRzviEVxSeEprGRud0ffiB/nlTdphTj9c5uQbCoScsIKqrORHXIsbjNZmmesel
LINdN+zWcoFZPQ9RTsN0lMs38tiS5nm9Pc2kB8rsLDxV3czoFpeXwPGfMnXezW/FHCPVA2LDQ80l
FJ3BZFzT1i00DIbrHvr8TWauQhBurYZoC7DlRQcGHAUNAQxcx6bek3XY1gzUlK8GnsGhWrwT1M4Y
EnnxoWnydCHWjKxljTAwMJc3BgR1tPUqLZsURUZMek3wBSvihlm2y/NkvAFL51CpA7vgqgZIbbii
hSG7hjGETJp7yvH9LZLQG+BatvZM7tpj5PGFR7A4dc2PxPUcyqPYO8uvt/teXtJN+WdFWWK8Uz4v
FMPRO8R3+gUAdUQnTNO/EYXv2TtnaW8XWJEptaQpcUUEcvKOt4YQjthHktYYgDy+BaKjH/3dxtiv
4LpE20BtvgtOwE9bt0KTbNOGw8QlY10KBO+4WtU1XYP6uuEX3568xwQ+7Tw9SZu7h4N+ZTU8xWbu
/QALHHviWk5RuBCLzR0JHEieEbJO472epLuCSDey3FKqQp0NckAWNSpMd/lfS6Q4S9fw9TySqxrt
FixTajfu1RQnv4msz/ycV+GcOIfR9pPdIYnT34rZkM1bdST7+Nil8/ejXOnrOFqIib21YW24Zmou
Eov2CkrDG5URcs5diKeUgh30JNDe5P1hr73oUDpsoI1a2YMiHtUwpaaKzANbY+tTBIi9TDI9ZWKK
97fOsSjpZ0d8fT+rOznhdgTxjrvm7Yx/0Jo9Mm0OadepZ9K3TfGbDt4ryI/leAbK/iA7gf/FFMdR
w/jxJzQxqHn7NMkdlWcFyXQhZHqRjukW8o16slL/N4SrHWcVeRZk3FgXQStRKDEWdGX92Y9vODCM
XgoBrbfeKXwxKwlym+Yh4UNGoi/s/zJDwsg/TggRaUJxKRMpDF5UJ8T3eaLDnWT8ux/SZQHsUwaf
6AzdbJtw5quYU2K1HDEPbnj7NouMErq9lRkS3z4p5HjtAl5oNdncfC0S+dphiLypVrS2TciMb2bT
Lm3VGgskXeuqW2eq+bE0cF+TTUvMYJ8cNi97mght39qKtS8oSN9lluK32VykUAvTmymyCS8wQHcA
7mmmCwO9UtqV1iVbjmUboa577tiOqaZaqpWy1yJonXqPxKE9Kz4tuuFgIYmnboIC0F7GK6n9DUB/
kxxmiCvxdCaIN8F6vF+M/Kdnbr7l+hE4nXy6fCJgmmWj+dq6qeGu48J9K9+M7PUXSgExojjYKy3B
w4BcrJPF6Hb7TMxNLTHM8iUP3ykphwhcdXlDuJfFIDgPuWVvDAZVBDWr4ysLF+7F3zmBF5tvw5Jw
zGuPcnMOaG001bt3Yk8KRF8VmFx5+LzBYym3EbZHTRXYHPMbw6pjqLGgWZwlGfGN7761yAYh6QMN
mJXj8afnCWtNh1mRPzz6y6od+a0h/9aKVm72OoGe4gq2UwefZ8M6xgLDvZKn83J9Oxw4bPpd9uju
fZRuUCjO8HYOQ4NVSczKmpt/AfcEOuTxLbgmcszVxZsXDsK6OojSmWXrODwGyQ1gIAbOyGEGPZPK
hsSNSvlgi8EZrWXoj/1JnqXTSacKvsFNVSVT2mu2W8iR8OKcgCSmZmt4NrHfc/+oi6sfZjs2d8dw
jKlqqnhZcuFo7xqVqHrgp1D967A+ZOWD/W1Doc1lalG8QR48+zh0uYcSFSizHz3/Hc0YA7n6b7UN
bUKY5GcyDN1GkljRABCowe2Thb/b6zdnkeoX+bJf6BEYgiuTgLjUaKOG59VeapcpU4zt32f+51+n
WxmFU+iNIWVRtebBJnCWjmZyrTQ4XMDfUXyQCXDtp+OJmP9ZzVedG3tSwoThrxyJXHoHz3jyRIZB
8DJma/45eWJWrM1qi0NtjTWIeQusMBp8CoU5PzKf3MJ/e0jatSJbudLVmKoPFISWfZ7+wf1eXBt6
Pr16bAPxNVUDoQmbMaCBazOf2xlZUcemczPht/trFRNCQof6rJz8trVMYPYvb4NlPRUJc4q6EonX
dRV3BfdwuVFhlPAuOvUiP44R3X1NsRcFy2c3reuRjThxMdF5WC8ylt91gF4CwAMyo8bubum7KHs5
OSrl9fMAV4EcrM3zhIA6w6VW2Z0+VCPU/9zMYXZGP8ovIuYBNaDxN0yMmge+7FInkrGbHTVZksER
OSw79/C/IjRJTu/ae5jFVnQygkVoiN9AohOJNpxn7zhXWxU+Mem7LtDEsmlHdoo5FpZlu26hRHLd
8BcO3fqN3w7+29GwfcFGze0ozmosg84MnWcgIGHCGATgJDP95Y5FiqfBi2CoP9vjcAshJLbByFm3
oyDPvCwsGsuRrG6ZcG+TVIreSdsOqXVLQlepGXl3Wj3wYQhgtsAjKINA9XVh8Jkq24AdMGIPZgcC
ddaQFTcEwaE/yFi/yn4q3r/dDLp7QjY7sDKyZht2FU0q/M2JHg+1hr8njEX9HHp6VqX/5riMFRTO
ZEwKeKUgbM5EGGCmOPuvUf7qVZQb2TrMDuq9KYeeNnU7RGGqhEYc7aPI/WP4ljenx7mCZlMLcRp3
X5s+hWjCCEQwON2+pDBWzVk3fXGwx8nTA92z2kalwzQhL9ra8CKPm11tpK1WLl8Cr3I/W9VqjXrd
BTt/7b8tG+2LHh6eje9rSGHvEhsQT84IOCZoQu06IuthHWyWiw1qRnUMoSOsIP6l5lRrc9MoXmDk
RamgaOy6gItjTk4tN6RCLy9mjGi8o0KwFJw54kXRBnLZJKDoyuK+Sp99DleJpH4upgx70dnngY3/
yIRgujXfc2P9/ZyhCfRlhza3A01MbW21LV5SIIROY+TZzoyVs2dHYRsLch2omcT3aRMQgEtu7l6z
DAeFGn16+2F9n7aaN0tuAWzqHovavP2vAptFra6wXIQ5bGMDNiInD0IHUTBeuPxDjWuamvNROwm/
HBC+wDiEGV7szD7065kGkHwIGsl8t9jShKxVFjIWdtPU9P+h5lLE3tAvVIifl4WqDhDrsV+JVkX1
Ymjv/G9/q7MxR8cIN6LJXwhy0Bn8ye55fmKQ3iKzDxWZMTIHoTbIkj2pnV7aFysrY3EvmEUpO+QZ
nPFHbMRukvLXli0lp5N5FntNVH/xBoKKRwvL8MQxhgbfFelwpBw4LSfCEoDQpNd8PTeZZZJz6RUi
jwOnI58Z12JQQ3OSSQ9n1N9f2wBG52FGoXkmASPWjD5FhfDEfdK5wvMjl+NHXWJ5zC/Y3n5sI9YB
WL0VF01UnrkpqyoXUApNpix4CPT4i5KZmJGp+d8aT2srgnFajj65laoVpiNVaKLIcnnrYw5wRYvL
SplGbSDGCLIKTmpJQySldur+HkRwvbB27z0lIsK1tV7aTnisX2v2B7NZ5iH46xM1tIn5VMB4/tWY
beFsRwqcnYF/BVnbTuJtWDeJLG1niXyiCdHISYQ8CPMm1VgAPueoWCF7OwXpUhKrkng1IRjL/79k
Hf95mE2TNFGNbn2uQBmXTLNSA3I4VlAHAOJlHVe9Fdi2lo3ArPwYeScb+Akk4JAdMDu0OSGWwlJO
SGgZiYvP/KbslKfdRjH27/KTUdTqyCCY0jPraIrchjhK6k2RyW3wNXvHzyQWB4SUrFz24KjvyxLS
6Qmhvz3jgnc3/6K3Ht/ycNmRrYNijwHBUcLDUSiKOf4OASXLFgB+YBJxRXtXY39FljdECFDcxkZ5
eMcnSZF8C9499PaNX7mhrfJv4yNroribJy6uEpoTnUrXKTa23qg/Qsoej337AYK+c8cytYjKvxc2
n43y8AmulbH/o+6KCHCoYSh0yIlxgG85UMIYkNU55OHdjuQuhsKI8pTuPJvhSmwvjDa3WGTejUih
lPQTa+2nbx822nDfiXch2XM3XT/T4C17q81Pvqp8GJ4ZP68+jLh6dx6t/YjagXI6MbNEA3gbbDsk
yayGC96EoZuSXhZM9JsPjk8pR2g6Ha6fDVBMu9h56Ozqct95OXqrwyC8lQrTNYXhCqeHSR1fxfs8
EHJs0Mh5+8JM6DSZif0VjnxUvwZ7Vi9UVyUA2KlUBamJSaeeQ8e6GoT13xDHvMBH6tZ1vuHXbN8J
H5PwDANA78z3FGaGbDXNjTmhtDMx/dPtxZ+FJwFZf1WIdbM1ZEDMRT9f9/S30UJoRlt5Kp5z3HC2
sOa8K1KvyFsREfr9JHmQYwzj8vfI8gdmwSkf6vRbLtG8bsNMUKakiC2g/5D+aYopWnaJ7mLNkDoG
EvwQDhDVk3bgTNfr+5w05Ti3Bk7E//1dRpq9v1DCEFeOqpmd4Et8ZBuW0cOz/O5/NNNOFnehZ8Lq
a37nxxald/3pzjM31znh64HJ7Neh8TekpYQgeZM3aucbfLucRxwgrJ9jTIVeJz5PaMqkpURadd1A
H83VZVqe6M7yikJRDZ313q4PC1k9u/7ZMhPZUMmbNHeeF/0VM5rBWHxLpcZh9rGzOEdQkxp1EW8m
YB2TjTX46OQHlMSciVoUv3cqWG2Hh4rpCUzJiPFtvpr7QpYGeN6IdqbJHOR961S8BNMLwHL4azFe
i5D0mgT4nOUwUv0a1nQtk0IUELG5oqNuBmivuZ4J/aN28Dy89nrU5Yi+JTfAWxntrhMHjIJXMGiB
5RzLliKQvwS2dqtVbo0A3vZgSN9NVACHsz5mgmZRnuYTcKCGhPV3GzeWT3UjJv2L+ApFzdwEmOdq
ON1z5D0gWaIfX9Uz39hewu68abOsw38zn9LR36DWTlOzpB9Klk6Zbnt2fnuZSRcU7KSAWrxprBgi
uSyMp6EXml3tFS7N3lNcurZxt+sUhjHNfkzjFytRYRfeNH8dFdjSKtmXS1XBgTA0crfOSl74DIH2
Q6SGHDO8Tlt6igYCuWyYmRzVa0SnfhPQnAYJFG1dOMRvj1/W8+dYtbzZMqbXi4VwA83BIx+rPT46
0PBvTknqoZpYryFtC2WBGstx/jL3BcYGOMzHfm4duihSG06Cwg7EoxA4WAJZicoCxrkyNo5Oapye
NvnpaEXczhjQwvz6cVgTpIkYcVpz+qBwSy7L2SCD0TCavH96F8YvnvIoZy6biaut6es90Nxptpsj
PVO6T79M3TSvEnRH/LSSICH4G6r4sGxVqZ+d0AlkKcFplrvhdWiH/ieO+BQ5yLgwAZ6hkOZ+iL7a
3ORTeMyZywY6bfwk+LfwF/M6OYDzmPYejqDv/JjaxUKxtVlbvZrgZRsuDRbLLi5nxMHLIvelc59f
8DJ/BoeLCoE0zMPp3xzSuqAEo8qXgIOXM31YWnZfOlXpmVsY0/MAWrNQP90qoJ47lLjyQ9UoTvis
8a2wkvmIcw9A3+vuOlHPx8LhCi0/cy4XIKVZOGTdFE8i2uCbZmN/8cnqeMTNu+yzB4u0gt9bUVUn
GZOhfLD8JLdmzEtmgUgTyOmRORBQCGrX4ISYu3fdMN9yw+05qz+pAuqeOCGNOLaCS3rv5BZSzsQs
n5ha6jMRpyDw5dnTEHJap6epRdPKOzAgzC3K5yGdjbBaKj9YqdaSwy6u+hIqmcUQUTUAstGjtAsz
L4rpOv9hINrY0plCYd86Ou6qb8XlyT7kMjjouSfVvFqJIG4AhovrdqRg3LuJim3ay5Ciho6HsN5W
MuLEb0p3mbfHDqvGks1QJmQXC5z0y0yXM2jp2IYBgFyR+1gtxwGHxu/QFQdeZs7zqKWcFTo+emCc
2Kggs5b3fpCihs/LNUZKy2A2emHfM4lmWsOlJQaBFUBn8hDuejBvhEg1QzDtWr+2niTDXYTDkl+f
VqeoOCRFJUFA70vy2akTReYVp9BVjmcM+CpORuzutWOCPB+lMgbwbXI1fpC+AzhuMwJAxQiq+Wv1
Dc8oOupP97D/7kg7W6YZr8+kyr3kb9EV77pBFkEMw1LVX0lvKJTMcxtlFdxwFErkb3RLpAzLeYKy
SSbO6+W8iHKSvAbKuyLuqxpqwIdPaxX78UptkggADJ3dOITH0R2wC6zaWMj3k1uzFg6TOsEGRzGe
pkX2ct1aiLCwc/ZPxyJncCnIwiWTSgoxAQSwYnMXkKRZSS/ldJrtsFg259Bpmf8VkcOLD7RM0WgT
5TjQY2PXNEyIQaUOxf9cwAOQIuWE/4TMDKbjvvi+E1QOLi5TsBcfSx8gdasyVldkuh5iLpa6Uptk
+noqYjN6H2ZpO5XJg+caRH6kdk6DRQsa2wIWea+msge5dtn08ANZoKY/n1EsYjf+Wgt0FWby79SB
TV6kN3y9bMDihQ3ATjeBQpdbOMoTYx2ALzVpkLhCOARDiw79cT9Syjl/ZBUdS/PMgw995Xuca9/K
eIsPv8AAhs4UdLS3XOUbpeUYbuNsaBCf1LZWMyPhdJqiGWOUFr41v+GYGszSosi0SvIS8laOjwXB
CNPRX/9V18Pr/UN9pUzxp/HeHFFh+xNLDQHbxFJVcGN43Crs2bPF1fItRgkgfVdS7feUNg1iCBZ6
96Oac4isdM25rhKi5FTT/deaaF0NTE6o2XOq/SOgYEJ5Jz2TklM23wXf7I3fupNjJRyilMNnc1JA
qvOxibMM7O8MF1CByj9y8QBFe1ID/5Z9CinhcLii2mVc7g5Fp5i/y9CPMNdDAv5v2Y0U9jt0A0Pf
P+8rhH7BL3BRd0liXYXETxlWtiM8b6hOAkDh0sV+UokRwz8NUMFv8zp1NgRDD5hy0tcSlJSBb9KC
FTS1T0vbIOPm4Y8iP+QGXxmlIkIsUz1ePwarGY9q6GFXwCqrBp9JE8BTMYs9Tk6yfEoQEFukgI5u
XQHcOyQ8EKcSpEWtHYKXMAnOGJvyAEc52XAs2LfvCrnTM4FsDTq3l+WdsN1w5Syme5m89XW+p8Rw
3cRnf8KNExqp6LixjOJGX3eV44g8tdkL/SrZry7sJjekzX+/Vkgs4b6/NTwTKOKZGhzP4vRxEbdi
6sG3QFo/N0CbuBEK1APUK/gMACXT0sRpl0ygbpMB2B8SjTQtIYP6UZkMv/SHiHpkUkSlkslqsiMY
g2zWzTeB5+DvrQOJe2w+EuTuOcpFHRbmUEjL0KKUwzpb3OrFiJzyBm+kn+FX25Cde9KJLAowv7/H
/ERqfG44fk/orXFMAykOn7FWdMX/mQYJzcRbj+F/oix8I7Hdq8uuicXwj2N5ECv/YIyppaPkKLjI
N61ioRwzDrb9Ty3CY0pF6AqKc2NxBU7v9svZkKRkKGDVDjraaGXCvt9+S3Jc5+EWestCYV6JnfGJ
FaZf+j39Z6MhTGzHxC6NePs5OnWTAo/GZ4kDGoZZk1aHVWIlvZ+SG/46tyz9H1Wr+0pjc6QwuOAd
WJagAST5UHfonpwrCTn8HfRYbZnMP3xN4zZfn6KZSyY1ATqH7nByVvxHLcYmDjRgckQS4LY+IOHP
Bl7QaTwMp1ePph5r6t3zLUhPAwjE4usHnCUJhW+gSLarTBTYBF+fOql+WF8LcoqwQ/paaIk7tPd0
hw8fQmSn8o7bpPslymK3ZUouue0zwPVVS3/vYUx2bSUkU3GBRXkBhraRM7kSiByXzZonyRktwDH4
UTOpQt3fVYChD7OhrHrlL4c062CElVbGaxYEScSBZfGJSXCrMDAG9OjlxDIDCJ4DTQWq0D44f1nu
eSwikbzu0iwsD+7AY+/+k0QmysMPS1zCHYk2/j2bO7Y7VUZxg/CSpqSKrSguSCPL/rH00vczRzcs
qDJqeLOvXytVVUuNEcAarDpCssRqUsix0CMh3K9bwyOgBoxsZFyUHa0NKp8YM5QvA4YHyIlHwWxF
CXDJisj2admtMhELzmzrJQ0JDaheLwrv62OeGkAYB3Sh81PHTfEDyFxCF/wzMa5c0vNi0BaOSFsC
Mg9Wlh0e6zOhtUzxjCXWf0aNIEY34BxWu4F4Ds1A5AcAnCHzntBoOt4HaBKdSKW5BJQFe2WPkG3h
66UPe2LJZD6uCq5Rx3ovJb6+LUJg3R7cWIhZbm5rZmzaYs8EyhZp89bVnowkeE1b9VwO0txKvCe6
E6FUL4ouSPXZctTMy0eggnRTlTYVQDT1h3XXKeeDRJrlcMs6y8w0xDVtr79LHZAvJmQbTCNZltOt
D45fXHl8pf1pi7/v/B/8Ar6I7moY2fRENl2yf1TwFyRLfKB9xc1X3kA+SX7ScEC6wYPlG52IiXsc
BuO1DXA378JTzQD2PsqtgQb/zlvYDgh+Xv2KPT3pPtaJPcuxnYzWf7dgFg+1+N3MSXAHzQ56nAxA
C/lh/YogXyClqBIqtYcgzooHng0VIa+vn4aulBZEZANqEU2lzpunVchFsUkEH6aNfvwwLv2mnmII
CE9Ma6fVX6EewdiUc9V85IAnP0APYnk/+bezRA1u7qoAfGqouxrwz6l/0V4gTvfrwnZc58PAgGXi
maBPPVyzc+9lrZVVlIGeLQWrbAKcZ552AZ12X+CpM4oBzbkSCVra6bbMI9IDDFsrp58oMj+aInTc
z69Jg9C/q1nmLUklJpnoKX0JTOfm3zlfopp6p/LhZqKh0YHwc9Dlcb5bmrmw30i6zyBXkKMBEOsL
ekBkDefZBL5+1Sie0e3aROymN4vpIl7m1ZdlcNf4otld+a3BLF+HRnFeAl8O7ThKRr9xl4kAk1DK
V34SKI53DnRJ3O36yB/21PZQhvWPpPo4UOngOZgtdU+R4MPWX4jZ13MGiodwhmcnpA041F2rvP8+
l1pTzNTps6nEgrCuIXXwmVuBqBmn2cMDDyrHaKVjR6v8LbRDWqD+YlThh4qEik+Yu6MoeP7RanoA
EBafKxAVlDjvZw1NlCMaOBET+wZc7j3RW9eOaaX8+oyY3spR1vdil0vwtppPnAhqcTX3PCQW3bWt
gx9EFazmtszzQYNHChKj4EPrAN/Jbhgg4tlxeXq/BFMRmGDFBZ3RvITs76Yek09hd0UrWQWk6OY0
i++eJlaCH9w3M7myfBaTQ84UPSE6UFPDzlB1ypfo/ljlL4cuHFotBhz6dkg6HaShhtyqbLNzVf6q
Sk0gsiXd7lzqjhs8PQr2zk9yahAMoMj5/gVOi9aEgt2r0SXPjXqJQnrjkdNzhVc6hBsVSiTyQGio
vwlS2R68U7RwIMN0WD9qnfgj39bSisGeHyWf0UCRsH9XvNGakdNboK2vyAUfVteTbvn0tGgzaAUM
P5uGFFZPUwoBBojYHOVoPIva/GYWShwfiCPUMorSQrLdK6Rsr2/bkWjDaRMI0ZJlltN8Kx2becBF
Kn1B5RcLEt9STxw4KzzQFKgrCfvwoMDaDTO+suhjtPZxrsYZ2Kqjvq4fJdc3+XJOC5AMjYFo6uzx
ADz9Vt3SIUgjTcrR+oGUvvare+bKVeLN+PMmLzFUq1w7IbI6cG2+DCA3G3ZMRpfPieQa9MAiNHEm
cQkN/aivT4thywTM9QP8amNCzXMRsIrJHqlpM60VAOEdrw/yW8uJT0ffv1IjLKRsl8j+ruTVN3l3
WfLLXgVmS74mao2TyOO4KUiJoLNlIq6kJIBLmA/Gl0V0GJCPifz0yVCAB4xJpfuDdBUvgUPX8dI8
UaXk0yo4rQp6ohL1toJMlWZxjNi74GFbRuGrPewFZ0IQA3dJv9E2V76ffo1tksDL9uyaSSPrALni
YUjQ3EONTxuQqypfDhlNks3Hq99PBLMCI3JfsmMgLKMyX6iYQLyWSOqov6kzDeDBCnM+mSoeumBg
ykwnNUYJ+2VVV9+gaWqyiK/9AN57+AMn3I+UZqngwPJuQUPY7msnEHCHvUJ38wmkA5GiFvRqzgwJ
PuHdj2ezF+W5yyGcpQpKw7G1Z2oB2b2n4VAkm4WPBJfNrvbgTlecRUHh3t6uBqWMmrCZ9MZ6Qhsi
1YvUVEsC+KdWPM4NCikHTWd/yvUIq/XlMRoV8Ey2zS0IE4Z6sSRoXly/oeE+g7sIND36Jh+tBWgD
M8dHPPQAt77yi0uf4K1zkz0MHngeXxqWUzOZJzdJFCM6hc7FQQwHMffygw7/dBMu+7ADg3g/r8mi
PRqXTCToNDj6fuHGn8ywHy4VW26xAdCtBGIi+6D1vWjgDmsndqraC8h8YkP/KvBDzLghrrr32V/r
14NsZT+JHi47wHjNbZ3cItutrqweelCLqrCcsLbVk/azZ9zV4pD4023iErMm08754Lu6LNnzOJFR
y00LVepeTydIzwc9kB9REsVLNKVaJuFfX8pDs20d9kQ2ZZZWbUSzNCmCSbdnVDjSsYdp7sNm0cfp
5mXh7Q3wIL18OI7p+BQiwsoUININgdWsPXWcHNCswJ1zg7v9EdyfOhxiQB7VTX4srjtPCxfTkB1H
wkioCne8Iq9nmJZ1q+jgAnRA3K6nhflGM7euNH/WjuZXm6aqhs3nfxSnmh6SY9nSLmYmTlOosGyR
+xAnQRnNtsJ9YmPHzmt+lX0apz659QEC5St4cmsWml4FvW0z0M1wCg7RmbEPO7o3gIguon3AHI+3
wyRP2R23RALBfvWsX5+v7PcMWJNu4vmgGcO5GtzAMeSih1wpRNYbnWcgVpk3eKqxMOjQBgy48DWH
FF+iknXxTOK4XifstgGSqobgxX/KyEMHVBsCzoEtZvc3TmHRMWczp1MN7LIv66scqIAIi4xXDnge
QVtp5JB0e4rtH5moPVMAoxp3bG/wSZOeXKJCGjT+8aPvQooR8I9SV8iNtLIaNdCWeak2PPuiSTEu
hcdMzLh7rX9+7ogAGt2gl5FgUTjIcgpZQD8t2q9lfjNQN4BotKDrakrNiIYLBe6HjleUFSkzhGNR
O5ZEhmaIzyfmwKTEThtp6bCT8SYYyFzyIqH4Kzs9HzCdq4Jvs4zi4ZFGi9VK6K2d8uxQ4OA/bybk
iIWmIVIfxI2EsHqwswawI+CL88JyjN6/ccRdx/3aPQFzvEByCMhh8JeEe74NcHb3YIs0uWKSDJZa
/Vc9twSQuwpPz6SIiUlKmhXzNJPIEi8F6XJlSnfyUd2Gq61S8jUUc1Z6YnZrzpDtRJj50owkbcoo
8xObckDjAHXbCHMRS2+dXyPUptGO406kihcCS9RpKXQ7SlUplWfLmS7Kg8UnHI6SpL2XxPC1S7Gh
qeUVfC6N4CYcJazd0P8HPaOxrcZY1W4IvfsUOEMdBSyquUiRw/Ys7M9TWGEqn4mL+AYM1+2L/WOo
GAFdYvEJWzLGNv2FS+9zTqqD4pRL11h2UGEEhoMLod13fRyDQoEJEjCN+2arkI5r5LB53cARow+C
jQJFoWrZvrcLS6f8Yt9b4RnYY4R97PNaeY3KYxk7P2yF5nud/lOymfXqyzwSVmonS6ciYaARrWhN
7CGeRAQmFxrgv1BWnWY4k0OnAe5gYDCTeO141UcErOiwiU68x/1Kv5LIY83wibjgQBE7R0UDFpRy
UerAZm2NmryprE0gd9XXOi/glWwZW2jepvynm+Je4WYiMTsljOr368fcW2+wftatd8jRj9eoPMe8
De05YtkroZLCZY4qredoF9c8Upt6+YI60cGVQo82UQBes0A8Qcqkz290bhpllDWCh5b34hFP+X3N
7VN/rdBJFHpjWw2l+tBMhhJt/7ABaJSuwUM/8QwRunh0tQ0H99y2YTXsHtvGSLU90Xv1Vbi/ofCz
8ok3XEjEncRg8JXJgmEuQkgfSBaqvZzG71onrogNb3p81WKyJEC8FyPqlAO/8tBRHw3y4Gf+SsTr
6Njcj0so+dy8SwZFPlyPr2tUf34UgzhKadGqQrJqwlnTV+nSkBrXfLYBy5dfbrax4gsYEL8cosxe
Iv9dpS4/ssVGDEqZ4ndPJ2GF15jbxWo/ElQwVmq3+RGOFORc+Y1A9cs/Kr+cjRHXYx7R/pSmOfXA
S+GX4n5OtRqUWj+FZRG5FzdYuCjRyYsaZtigblyK5W9/WEfNph0SDX6KfhvYSwseodxI7iCUn1k4
NjRYSKbpH28uCS4SrCsAYMoN5ZHb3WnhJVbOgLmcypIkMBCk3OiKq8VUVGa1+Ee3AJRPFYkJem0o
EvUgxwSqC6zc3+1nHDNa0fJlEfLdcwTNQphhpgLquhbfuU6zmJWKQck6P6rHnPWsPda7oecuP9NC
PXbkg3ro7cAiVnHwyN2IDmmhoFl4YYlVZVIYPwd//vTI5eu7VT/XlEVflBlpNIGghayeE5rUQZDA
aa+AtkJ2rqpcPtFzZWJQhkQR040QBbq3W2gLpGihJSg0w2PzoyxZv3GBwodncV67x3NKUGH4c3Va
SjxFhwfzA7CISBplc8o4tK3u5qn9YZ+rpPCEZ+GqCoc6ess1YJxBB96xaoCZrrLXhcNkcIlTBSin
Uhe61gWhc8XbBIdpart2IcSVDHzfSJ/2OQMTK9XNYGRow04S+VwSO5g4fZcckU3cvCCtkcYH6qIa
Qd09kD1IuBnfP8DiTTXpPpsO9whzKJAyDpeV/jtKYz0gPE9tIfX9dQSz/SKS5iFQ62bNa7NRhBlr
A+JKHTVRTz7U8Tqay8wNorCU3ZixWEZKqRuYSlhlJNRsRiydvXDkbiHGB0B78iiT9KtwLph81uEQ
jILIxf+ut7YrYF4u5kuazqPIAmenpmGM5iPlOeF71hIfhoaM2Stfdf3VqPVk1Fke1/tPdp2bX6aI
rvEpmmVvtPyrNWbGvyIbu5Uzi9ZtFE2MQL6hJ5qYgAwyuKNP9g8UpXRIeI6TPVtwqztGoPzavTP4
VKekHPKdccLLuT7LNJ/snO6u9uCwc5TUSok3FmHo54PpkZAw6PoOwVEdgmd0Dk6xQ+4+eJP384XC
oWuDuW4hF6Pg+SzvxI3BPuHi5smMbgPouvwAma43F5+zza/xezPYPAmaZ9O6fATRAm7uviPItNuP
HcV1dwFvPeGhAyhRxHcu/SG//62MzRkR1Cgxk/J+7eKE8dvlaoGM9wP9meFGT3L1yrROrQLWOFZA
ZPGV6FDkReoqj/6P76oWsSdm2et2vLH7HHL4IJLTTpnYe5eRlnHQaxKh0nY0yn5KS3/0ijb2bTv+
ZYR3s4mxsgVzhJEymoviFDCd1dzaCnjN0UadNqQi4rByALKHkao8sxy/FQ2K5476fyDWtxkQNmDk
BQj0jzjPj34yWTRKE6atVwMYo1MyqKQdzucI8tENJ4s7n7wZNFdavsJUUpjlWO9Ya30M4YqA/X0p
IYrqo8VZVaKXtc0WeRXtCL08gi5IqaoXsPvP6y2C5uUSRWa3oDOJvRev65ezjRq8nKZFQmEpa9gL
gwvUOssaGt/o7EAWX4uSuBovyrUBKvMwO7xhhFSX973Iv2W1h0lAPN/hrFHc5J6MBoRmWlv7zSKr
RvYsFmIsxDIeRcar4zjhHG3DJB430jVRMoYOytfsUGoD3oa+Ui2jdEj8a9ng4kVzA5rToi7eRES3
U+bLBFccZLOrO7CePjox+xg9i9iA9nBhALTFy96b2S6fUKxPXNfq+YQ6NJ7Q0Kokt4FXW37c2BpQ
+WevxZ2nXJyxaaAvqlOmrekf44P7/NpTsXUtAnMR3gG6IF/oGTrjJ49u5jDHCuMz0DPLxb/2KleJ
pMUQZNvRnlUBbUCrPan4EXCgmrp7NRRg+b5QO1vNxbBtHLCzqTKFr/GGOtcnWc3uUJatdHJhfYAr
pVcxrjmKDsEGb4t53MSfkdjYwiRnW0UiZFqIL3ghDwMOExE4lmYnvzTOeQfd3WSD6xqO1xlEcX7y
GCtkgNbMmBtnDF6z5ZOEmzSHwbIw+k3jlopun4Frd4xIPfMRZzoqoQtvUtBYu6KXIWgH9mqokuGB
VaPG/6QNkh855u5hQDAy+7dMhWfWOjuo1L91EkXDiePggdzYM4L2ySs5aGsbG+kxgwN0EsWPWJ8x
Hr54rA9VOAW6j2BX3SFfn6UY/P0qF2Rstj338WNBQEvDtIIeDxjKSHPuDwhq4eMWlwFFCbolT8TU
KIJHTuX4KHsHF1ikET+nctKVWCd4gK4Sr0dQ3KpDycWYa8G2cgN3RZP9g3uK2j2mvXSkzlKRoTQz
eJG+oKrX8Qwq4to15in5XoLI7EKzxASGMuAlf+60uxEMvoYqr6bS9mNzQUfZQ9gRWmV60hMyTdeA
WlH1as3IbEq5XZpvakBdJgaeHtZDKihw19gcmN1QxF7f7qMvxkNhR0RTo4EZ+x8jwPrQhRYXuSfp
/vRokK9NfIJNAHZUATGdRVAZC5bSy2ZvwmGvmKq3F10pzcekGHD9jK9fef6iYT0TYPfWuDMTGZ1m
KqzTvu3VIvsvqKSyKCfeFmdIm3cM3z7ljcd437otwzuMUkitkCa4Zib/Qil6U9yl5xWvU3ftQP9t
yozYl9YwJ1x/I77KittpPmTuFMsX9Do6bBcafV2yqsKTgunMHt02ZMMYBCLmPffCg3HHBOundMuW
2jPAY9dSF38skIm2lCY+Y43viKZHlCzjXlFneK41SqwE075+fkwAWWs/cFY0ptVcW9fZ5UatX2wc
9i1Vbzhvc1QhJTLAaFdgX/ZbudN0hRFHYvnDqStxJhZQnQ4Gwzf1RvHq51+WwOC491MVr/rqMbpf
SuIxL9Ae1gB7dlFw55NGMbibMqcsDAFJpSWUY97w2t12CYYbRHS07SU5IMromN6/wgkk50fo+/Nv
a2BjA0TelOMCZ98Uwq+NkyS7H9nVV7B7fD8OjzRbWuP41t+sIofnT9IsLpgEKvfHhwJWbT6wmDD+
j/NgPhjQjIHDDTUr2DCuweX9BqaFZUkbejCMdf9hJThMzHSPufdwo9ZgX1SrtPViL56xqkjhizVQ
KGHil+0mmO7Pzyp3CVJ46BARKhO3IrdVKl1sMQnD5gOCLEAJJTPtRF6FxHOAGL1vBLAuXNb15jdA
VLcmcG80bgSab3khW2FGtBcNjXMvk1rD+1M79MwyhYyjh5dHsonXqWceQqU4ff7jpEVgraWW4oLr
tLTFQTzJer28FvQRi3vRtXAlcUlveU+uD+kxHmzQkfZ2rURE37Gu8B41DMAoP6b9GMqmDxQDqOx6
6lOLhOHLcZQ64b0fPBZq97Z8qabJb37mVnf5/VQhIMsiWVljFAK4h4efT/hS6nhVim8bEWj2/equ
piAPe5Cfubnxe1V1snDSgPmtt5U4VxFyV/HL34x8VrwRQwgQx7GOZo6PuU/yUBDpGFBnKiLO/kEX
9hfdZ/Ad9vojLVe4HlbZnIx69TXLBJTgk65hiP05W2wBrNWjKKxA9EcyzX2oT/AuaSIPTYnCOuGR
HE/7+EQoQkeWbNDj4b0EFNzGIAe2TVnJ22hNwMa/szgUlZuyIxOECDwrHOvNIJUPQUL/2Uows3n6
ZfhpyC2/kv0lcGRyK4CkfNx2qnsQe8MwL9ePeX7yZre8ZYPQuv9or9FW8m2+JZE2E4w2qCOsldAX
V875HfFLNU20oBexXjs/iX0smScKMX5n6ZZY6lWhIRcVjYh8sEsgg1vPvw9qW4S2+iyRyHxkAlbH
T3QpmQhIckR3AItvecz4jWkuTm+8x/pDBSxndqRk0G/GD+29z7dL6BJikGy3prd+o7iGprEtH5jg
vZ+5/xYXVFwmEn8dm8+53EDuHeaHJy/WVFZ9cx26Bzq0QLFHaamalYh9zbYVUrZdYLW7tdnL65XN
iYvhNkYcQIRsNWTzyWKFYTS4iKFoLadI8WjnvP6nAbMjZxlihoBB69Ggw2g2m9+pDHSpUNjHQxNs
XySlWrC0XXJVEfEvfoFS5S7m5GqIB7e7q7jeJXZOjt/4FbuMnfSogZ7/bGybjTqgz0IaBCe/jJ7B
aSmBYFmpoPIBRrtCt1YYQrLIpxX+YnD+waX+Z4kbltT1nRSwHug4J0+kRu3qoHJYxip/rozaeQhR
3uFc7/MT0O7O/l64LT4gRZXgzlmk1qXDUe39IZ2/jxabVTeFoNqEgaOHww2xP6Q0VOEY5+NJEBne
16H3ZNmKGHwjWGEvpWdMvhYF/jE56OGcYDhsqlNT0CR7AnZzkxhosyC2eGP7KJF3D3lYt3usrneJ
UrVP5s3yVAHVQ3ZQGGAql1dteWVR3+2e4OWuXASPbAYVO0OXggvBsKM3nQF+QBs+UwUZCqJnBwyX
VSMOt88U9Gy14K2/WHL2HzU5t2eCkV/CVc6kV1gPcKJNAcVSqgp9mkl9jR/8UZ4iYCN8PxL6PUuO
UpsnsRPbxs4IlM1DeU8PcBFJU44Hv9BbK0h1jyOBTzdSMwWuK4rrc9svwZ6GHjs+ErHZnRvj9kue
Wgu1AwK/nKoe1zIB/FIr/jSESLbjK3U4rcl9+bCD0cJvs3FzsebCbUT65lXz4BugQcAX1ZFSTg5S
5CS1eIZMaeFUZfqJKHsKAMmYbbk9wlXDmnagu9H2/uJBTUw0KB9QeaYUrMYNrs+xgSY54E6qrKTr
8rK4i0oyml+pXLASZAX5IDqvHOpHzoQm3+7m8uW3kZSkZcQHlmq+BzHZA+iDl4G0eCxW0MtaT6Zg
PmtAcPJ8Zxrpq2WfjGrYsslnwXWxPar+YZN1elqKgxVWKMBatvo1jjtFBO1+QLAy9AaoHssZoIoh
p8KFsQRJKnT3aJkYSNVomEHJx+cZ+NIBiPEPp+EBPDU/xAonfHpS5e7oX3pXVEpq6hLjf0ULxcCx
nuwAFBWx1+2tLFaQf6Jratsf+574IXiunC6ZxfIR7s45qX9+VWILpawWhYvYS9GNlwUulFO44ECz
koOqL64GFyQfYeo2wG6BGZmod07hmTWrUXvPCtNrpVkjFwveDjbB8yup3QTnA2qqkNw5bnirUCJE
enRDI8lfX/NyQ1Mg9WKvNDB1VM06v5XOnQNTFEnWqYccNQ/MZFRtOBkWK47qcJXrEWXbSD2uQ7WO
XTAeCytshnupjaM8t3bPjndPXQxaVqVdBP+PsMSak7FvxKuJj5ehi69OBU0rqvHbnDRQOZCcqlSS
84FyZBovuWYeaDbofXpY2yOZzIUzu48y/lVRosbcML+fc1QxlfxyAy3duJEiq42oeicvuoiBhngd
GCzbsmR0QJRAEMuGV8AqtyhLEuxsvVNg2UOH0IN88svAtOU4LCI5knR2n1ZFmIc8hWaGmvMP0KFF
ER3i5ITgMSv4qsWV6Bu0WmyP257VF2cAgrx3A7AzqfXd1HdcH8fgXbBCrGDkNEz48DCGkbLmgYj7
yysSBCici2lZn/kulSDO+1wLx1V/PCtVYe0wukWsp51h9/jzfq9U12YP402PsxN9HHzt5iaOizct
qEfXCHCzy1wR8nbrBi1/ZF5G3BzAIfPJSq1OVDsjQcsJ1ygU0KegsBPwxhYCzaXzdDDnjvpcAO9r
NRc2P8JjNdwzDXkJKp2fn43+96aTDQNuL0GOiYTCgFPNaT8E2qmjjbDH4mSdG4vu6j4dqITPJgJP
lZsHqb+Xo20RfEbml9gGbNu5sxa9yWq5pESgQ3LH+bH4F8qbZH/YErweD+wmCeuKwO6GJeCcUD6W
aSMrFGVIaGaKdfXeLtFe81s5EVj6drgluv9aXuJsiwmssYt99vj/1TDNbiCCh410J81zfUpGs+ZL
v/mqJ2ys97LdZ+Jr1mih+Gf67fOD4XX+vICrx4kjJufHCNCjPXD11CC/meKJ69HmLLlVTR0Kmigj
7QV5KeSu9gm8KdOSZjn1Ho1Sg01uzACyD92K/0iPFIneKo9+V2Acx08D5xLCNqgqjdZsXe+3BWg5
M3w/+FzcyFd0yCQ/NxXbEmLoPeeB3apWan39aZBiZNJ9sDJtoM2GdDp4z5BM4du9nqXVwBlhM5ha
3EjtPzFBWm3gPx4BIHiVzxRbHXoF830BBrKwX9gLIUA14bFol6GEd6ijzCTY9EZUvqI1/TfxoVN1
lcyFOQT3lCAid2P4s4sbGp8hSlRmktvl8kPjkZCfPqDSKvb3NcJYKvQIe+23H+KlM+d/Lc8t4hNG
JrBcD24ELQpi6iJAbA5dNyIx+HKLAewgRUDe2Ntp0egkQ8nI8u9XrX1UE52jidPZ0yNQ50PppxI7
qrkIyJEQ2Z5o6looXVZC/L/OIcMH38yDMkYqQ+kYsqv9NHhXE5Kgiun83PPkPgSwTihkQkPkVM7P
QQyvehuCteFAqAjb1r0ILDpwJDdNsnvwC5Mn1/gSggUaU3BrA8oFQxcktt9/hjBirgJ0VtEqHX5D
37K1c8qPgHi5CO5+kU4YKgCGlv7dRqAY4ITVPJgiA3YNFFMZn2KqDLCW/pYAjKSzEo3C2wp/qzg0
QwTypf4inNlP405ndP4kjjbphtiJ3HmsiHYWcfmI53DRKqj/ULPSwM2ksoQAM5cQ2fi0ZBM6Z4kp
xH85iud20j0JVGcHBhF3Gc+WriN6UmnQNL0bCm8t6awF7z3CrOiuWrXrSKK/ZY9WC25v69YxjYA2
bUMnnRleoIAo7WeMJ82PvC5xmBRzKf1aTuzXx3AB+g1HCxQSLf+cldmft5O9WYZ2nBLkJzvVp0kc
IgXA1WKT7/fd9QxzroUjFFrY6xJcMYTk7DChO7il3XGzdBJ6Hyt6tiBuenBrcTyzbhvWIbIyYlD1
2FePbf0YflWy0L5HzKjKpyqAix3CsAG+gPHmRFsBKuGS3vyG9VcY9yE7S/nJ4cjMAqVST+vW/8lR
2Ccxk4fwRlrQBdqPM9kKFOp1lJ5LmIrK25Utc0lDqy89hd1ZJjV7cs9kkeo7suW69iDw0EMnijS2
K34rzTYOv2RRs97vebdrRLUUvYOD/7wp798YXJLtOfGr7iacjTHhhfjf9Y8bD4clL62n7OWIJXoZ
1IpPE6+ZYlypw+jOx499qMDoZ2G5x5/MdyhBW7S1B/7KhocFYTuJBNcyp/HWEpZOKKPSv7qAfGRu
DMV3d5rqX+qqKknHo1wz1ny/GU9rMhctMHUVhryoqNmxTc5kpHuCZx5FHMVsqndCTX76zH7pp7QF
sqmbIAIGJNKKJ6qf2E97YsyBLbUcZaNveFjhzsRXI8P5rAsXIB3npekMXyBRJYFF+khhh1dZn13U
w81I8oVx7qGmLGUr0hCAUgBV+XrgEhY9BwtCxRCOdNCINa3H0mv4aox+bIrxQ2ntVIFUCDPY/rUR
Rvf9V8Y1TakyyPRUsrKnalTFeHhxSkD0tw2B+FprPWYw/sbhQBU1VOSniIoZcPA5rCsGJJDG0qn0
k13QueETP7fzJ9NmGuCvms+k5QWD+QiCsAJNLoGETBhjYtPl5wXLpGSmebi5ZYaaV6vDt2aJyrSb
egPSLpTuUVOBXBS073uLLFV2Y5MzRSako3a1/ZrCDLSAJmYPgFrVq1t5X0tOAWafB+GjELyVlp8b
/6SfJ1RnP6aDVnWNnxYyt268zNHVS6cj+2Mc8sRqR02tlP8gTNBL4H9mqzOpl2plnEkDSb7oaahp
TcuPLbBTyTLU3xL/bFC55U8uOgZmgw5r6w2s6JAmjGf/bzkImtVayC1qfRPxRgy07LnkztIvzaJM
UoJ9YPWxforwSerfxsoTd0CfH3tvo1VPiFL9cH3TD94TG3V4dC+BkDD2qgcV4qNbZ43A6eCnQTc3
s5kfyZfI6ZhbsroiXuC510wU+8dGklf3vSnDz2RX6PJP95J601d/8dQ69a3cHsDVVJrzWcBM+qIh
BU99j7SYkLnZ5o9zqYTHSnJJ2HS0KcH7v033pWls/0yOpVuBiLTHJ+ad9BxzAX8u9RuJK8Z93P6+
pcklwPAEri4iY/SoXdWKU4f6WytOnI1YVDvulhFhZR8U216tIG019sL//Vm8ZU5XmmWYrHljndjM
wEzZ7cB1Ap2iTUU+IB9HQL/m+R4/50EgLIBWQ8Hyz8NAJAR/3LmOa/JGlsyGGI3hOUUxSlnKw13g
fzSETsOUP8YKpVZ+lu7ARzcSpgiFVzTFAmmWNTSPWaTf47m7E931TAOTCK0pW/5b8NG9fg+klmXf
6YyqZioMN/UOvkwsf2z8ZjcgXU7QTPpQ0WfuGe7A7ybbnMgz0tL8hfRiwZgsgd8OnCG4e/Y7L9AY
TYFMqwVMR4FtKDpaLrBnR8PdfKXsSoVnWqq79LFHZz5iKKJMFLW8INfcI2n/XlLuxh4cGEJlQyEF
R0uqEZyBq4Ahu6W2ZfQBgMf9F+Ovg7Tn68u5xQ6DdInK8see3o+UR7L48/zrBtj/kWRQ/VFwzIod
sV/HWiR5H/9LvmLdNakzX3Dt/a6hZbyuPxlEGQ3VrurctgbQUiR1RVQXlzVnOar8/mbG02p5fMn2
wV1J1plFwjwaCQJTjBRw89jRdiX487s1reYebyuNIiRLCY4DxkckRrh+qTD86NvM7putMmNFoUDH
PrXr+MhGWfpSOcMiO3CvWo/YG7Em2Nu23lV1JxoZXO/AnaUIzqZCnt6E5CP7KYn36WDOTkP+5xpJ
36nYeWHBpcXvikz6ZVxxV95hCWb64dN2TPd2cB566kNTeOU8BEDi5K/z/6D3NT0m8TouPYiLwZmD
PSpiKnpz3jGlkG4tzqFCrBFqDqBnjLy/wwZO2I4Debv/NbcW2Gk+UAqlOlBXiJD+G3Q8Bc7j/Tkj
8XR+p3GAuHjYwbcXEQCRJmCwxMHb5ynymPgw0z/9qNL1SKgnseh/rhC1HGXX9ZLx66a0BMd9r2wT
3Lm1vfWOnDBvGmEL4vXrjE51K+6uOmKacqcaYi4iLZNE185OUVgNfrTNuEcc8YbpthtTU0z2jjkc
1cl03Z954nwcRycjGHl32HJdRt2sE4go3UUwnIw2RckqUdUEQI4ASqQBJn1NtckR7jWl7CtVuO0b
GerMxE8nd5RS8WRGkGzf9qgpd0+yzYi/N/BNP8x6KqdlhrIbkCVkwena3vJPRwi3sd5/0XQNCYh3
0WZvru/aP2D4iunDqDx0ynZVbMjEz29YvBAXbxrQKRjduxDS3UiVujX4uycMprqPLzLouRfDYoZX
ra8VGrxIAShC5v6XnJ4Tk1qH3QRzTj8vDJa1lh0wwiRabJqvGHUixjQv4SAcohxLUFvb6rJFaLIm
T0Z+s/HetLQhsSwZNO2q+w+IIufhNRXQQzxZ2b3I+hT+ZPxhi15CwR1RdpagTH7nkoeNW53OV6Lu
+slIcebwcCZmg9bFNJr/72pETaU6MzUH8caFpIv/PY8LaeBAzdQIbyHSP8u+masAfRTLglmYenIa
GCHW+gfCWtG4/IImH5gHKdIvhFv4+QxZgaaEP4xVLmpA8TAM9+LRv/tydOgHuzc/gP+vurH3suxY
SMflUunGqduqmdZlpKrzleysW9Zr+zVTezZMtuO9hMe6I3dcz0yRCVN7QLBIV17ZeEgapwbR7rmo
Is/PZZhkjP8wXRp1TLr/I2kBt1Q9xh0AD+fS1burywOQNO085f25gFkQe5/KWCkPpYFz37zsxXy4
bA7q87tfuNH/BMJ7UTBram5tZ0PdolXrXvMi4scYnGpsYTEEDPD1IMMacX0dndi+dpibvLb0lU03
QiHT//ELMa8iBzV3pEVUerHkOQ8mG1fywz12ltf6fLHyrVYhePDVWolqD9lVvvywrEFMq+l4khsy
YQGrP7KKPI7iIjSdb+yMVEh+ABiLSUPfLyGaIk7jt9bVvBWs5XOeoLkxl67bVFKV4e+c1ZzD1gpu
z4LlIH+zYhLWhkMBTVYuNOUtOXVz1hrgWrFTpsHWFIa2e4ZB+4R2M3jQW3FKve8W7gTsnrsTrViE
iMTdWIWrKIBpM+jGo9L14crsrZs9DkYM4bzNQMxTAnKEi+bqeRQSvieK/8tLM6e3Q3qXF4baRkvv
LT9PnOS61aBoezLcLdxz9/yUoBgTd/FMlg2/mbzL6gyYCNAOmC+hVgIGQ3idQHelwdAV70H0mlEW
9O1/C5ypV6uXHDNEOZoFhbq+lS4D/Pl8ZjPMG6DtFJJ8ECVYR7+CLfu1YLO5W7mwjouupmdBduUf
XLYK0A6EITNevhJqLPMzN0xJRiWf6QbW0TvnXc3jLtZUkvkONQxDPkGTMLdqMbciPYCvcIVgoVpN
CpNrUOJO1mnOPzU9DN/6P1HSHSbKfcxBCEnIehFBl3CN0H4zyoeOCW8VeBsMSOS9r5tNtnPoJS0/
XI40L8AyRqw+i2i6UDrBirFDcz0nK0IZYyC1Dabjbmi0zDNvb3f/ASclVFt4AHXH/V7z9ujyNvUx
IK0HU2HASLrD7/7DVjuoAs1GP3tO/ctrNfExdhejYqiIG3ISOXkxt0bsLbEjIRJ6lEVfVzM33Tac
WPZb7rp7QD52aIMoWdfhPH/9cyXDEuFV1nOyrdV5OF9M2LP3hgoWmb5VEBnjwbxOxb3P/KSTeZL1
Sy0pBKHqhLfUeSLJC4I0vj4jsC99hChIsx/zhHbg2bKV/ILvpLElPZAfbrGcHt+HeawU0f3C1Kui
FTWV/JZw88alYk4P771AcdEblOFAuQEtOQTxeWFBz2kcm3SU3YuUKh3PTzWjyUGJUcp2j1x0h60Z
C4lx+HQmcQyFj/YmGzjI4up+uAouRgAYMW8yqfpZlPYYRCz7NZDrYjHsLrPbbDY4xvACdoE6HS6Q
1nGgBA8eekmMNE9ZsxZrwkBRdsA+IMISESyotnZ+x77rGszU+8zGNeoPjBPcTK5CLMdTMl+iLhTk
k35FtkFfEUfbjYKTSrQ/X9SmYUznSdwRglgMUe2ji9eualUcDVLxzz3nQLMFsqesHpn0qFLt8S4z
Xmsbnvx97qdsRsySXFJIlQncYVIZ6QKl0Okh3ThfSgmhaOpH3UnkWC8Cy1l1ubfX2hlOEta/DCOa
zk35TT8YnV5ne1kW8Xue/oawewBtm2EZdJhKLvfVqudqsdyz5wGRk9FFgkMwHPFeUnR+EMp5tnpt
XsVxWmAmGMA556xe+14nvpN7YFAKBDqvlNkGNIwvtZPfNFCXoC9we/pO8ipNvOwddJrtfLCxbT0H
k0IqH2akCXLDD2Feg0Z2JQgjidJgwbuy/NHaKsgVqCPT4NOif/inXcIqUqsIwf6ZqOvzhoUHF4qs
TnxIIFCsV4xA4lHgKmKoA4zwvMTPJsnMjzBh6svxgbJOAIEnixn1jfgsHD0bTNid6WJkqJMKo6tB
+ho4os79YgZeSpoY5zPmtU8DXMWAXR6pfFKJRLum0XVyX14N0xHGIgXw0CoQzGVw5uQJFDzDmkPq
sOm9jv6HquI1UVZi58ODfpcNz2TKYrfPMZquspAQCQdMaiD79JR3GHYHd4o/HlbmbfoelBBlpJ+O
XQuXAN2IGW9za+rqnALHt44CkJedsJdFukcr2dNUzs3aubtwa6hFHDq2RJzvB+00Vsb3o6tZxXj6
JliF7ZOng+KzaWTbLuOVf5V1+/F4/JtgB1mZqEZTwFqWKLJaV+6VtLzXZYJQ8fcZ47jmCgP+KItT
FJrI16pYYlb9Vwbiw00S5GOgvWVZJQoEd50/p5u58Ri5Ohr8Sdl+O5y4wQifomMyEgKKjMwH/04w
WZ9FgLCQy1h2dk5EzPSD1PmU+E9cjW9KiltNyuMCrijadw8ssc/plOoE3n5t0RuNeJtN3ASNfXxB
nFEbyGTjy/PvbK4JpxACuTgEv3BVxDaUZnV5NEY4QDb8Yt2q/TdBPMj9YUKc23+i8YpGliBUIwFm
wS8GNZcoVVfO6XmdD0H4MYrxPwRaBgJnZy882iyRkM8mnFXhW7yg0hpeuMAMMJlGAgCYnqPisrYC
H3mRUvLQdLCpYXauT1jdoU5D2gny166o+yrEKJ3jHCLjhO4aH89pSpXJ+e2kKpL8YP2cuDrVXqH3
3HpBuzf3plq3MhjUH4yPhyg1zJOYbQxlZAtIVNcm0ZtuO9lWxzo0Ml9PFEEI8BQqQ+qiWM3wCwUj
3JdLZrvzWWu7PNyG/5InSMJP4zlpIJk/BWTutXOeg3treAj8t4humEpkSTwM4H4JObfayniN4ewm
I8PPb92Rr7RUmq63uo1brqIDVvFKKYmZTZYTxJgSAYaJ7e4o3nVLE7XAXqrigWWZw8Jk26zRhCaj
BFvpQnEZQb4IY1r/5+wnSeT1KODu//xoLgYmNQd60YFWHpJXhisvqBu8iyjyQhl7vwmXQzu/z4a5
ILQ3FzxmINzB3EJwr30TkZAnKIdS6M6AJMsD1miIGV8eflDZopIbqID5Rexr2ZcYhVl2kTyPa5wO
WK9tem4dGrg/a/a+esCZJowxyEssK954RyIVut0nKw1czjSKWcYZ9Xe+rGgZsygzBJF/86XKL9UJ
MoOuS20VbFw8uUDMfU28DeG/AOWv690N1t2/QTtc06wJ7tXPm0o/6CsHl9CEXE04wexUpcEW6d39
Ljez/i1UsK7Q3pk/4933XJoQXSEMIBSyOjcw44YRhcS2EubGpx44UN86fn/OVP4bDTq3YgvtMxBM
178P+nOBZZx69ln+hGNR9C4htfWgXiVcoJTkVilrJjHEcR5MZLAdcy+phmQ8s+nHQOuMtAi+tdFg
5VnlYCimn1aF93vXqOSCX36Phj7l/+zGwjrXcQmkEkXhRkI3cTz4GMX8xLUm3k22lCmvNAhCr27P
WC/LbBOmo3875cWEpUJ0SzoHXZ02s7XHpISBBA4ftudJ5ZwxkUW3/Fl0jqUMiPM+B+qXP8+Ki2Vh
lQJYudkPWxrsjkyvRD7n2Le5FZ1thvxpfJTv4Fm6JJ2erBC0DmNCexMLs8ChXtPaqdZNUD6CHNpA
Xd17AWrcBTgSXFKPsnJt0R9DYJt1rz9FVfgTMc4QO586iloPqhz33FPEvf5SoneyWUgUQJHzeFxr
Ye2ZWSKx+Jh6d2WoGzdlf+rcdPmrRPNJLYb7xYIJ0jPzbBSPLLJACDz6UewtkZPaIJhQDJFPTyui
VgMNrYnb1hilINVw0UUcoVXVSu/45N2XVxx9O9DByb7Av+KT70kASjvyANZaBmAqmKDubx7uzKtj
0z9kLutW1KEMTKt2lYKvwQfDdwnw8z9EoaZdokUY/7bCNafled3SGRMn8vMSIyth8ZFWgfAW6dty
zyEYiqU9d8t8ClsdRm++7oAkGy2UzKxhHnDc/3a+KB2Lm9yuQG8EQutlUnjMjncoVk5BgP8JcpTW
SE/Dv44bFd/QOQg0Nms0bOvmE+tz0YhObDmr2BWAh1/unsnJPsfrVaW/sbVNktxkYmCqgsJMgjNx
qJ8x9ZYsOoO9AxVQNOhHcsBUJsXoocD8t/yCHK2wle6M2WBfGH9HQGH18PXE+plHkm44OW8Rr2zd
A8mwB2ClmNvfdwA8gUE3lmKFcER6wg6DSriFStnMoeX+8nrumpJP/vTHE9NUtKhkTXcH/wDggVvi
TPout57S83f76Jk7RNv3nW0f/F0eyogYmWR6yOqA8BpXEZzPG5XGpRAfClehG/KM8yMMtOTlRfDh
ZoGnj4ExXXFSE9yvSLlnaVZXj/dB3WjkeFH+Nctrkw4f/6baw9LcotnsMI7Yja8lIZDn2NBQ1BuN
8y48EvIhTDcAVkRb1aO0tlpJYsRWylV1KQ/8N75GCDMpgVDZ8l0+gC7AVv4pCFUAVz5X36kED4SH
cMhw5520X0jD3MUJNngU5cWL+8B86IW5RUMLH752Rta5wIz0Q9jUHnjnU6E6Re1XFrDFWcqwOerw
0jdnpOGlGrjlrQzXEUWGvF2Y6svqWfMFqhbbK6YMFpNgqAqWQAMzC0QUjqUvLwxDLmIEKbmyuRYW
TlDF04VB5NuuAIH2rk25eSWEZd/L4IsaoTFnJQ+pmM3e+pZ8JAnjQWmqs62SRD2PSHyRNPhzcI2f
3ObPd7QZRChlbJJhDGkozZqJR5WQjjrDxTp7H+Wttdc5zfdaDVIBtnCLlpjXxxZBlNqBhqM0LZ9C
j8h14qApiYyt9lpABwbyR4eYe5kpyQwOFZWqrUI11csq6HRU3GbOOKRCiFAz4wOvXZlC2tYq7T9W
cw279fHuCpVSIOs1CvvJWLipH1S1jVn+xFfJk9F/p7A3dtG4Oqfp2bpAHSU0bpE9TPNL4YLC4IUZ
jQO49Wi38bV/23C9/JTKhkgI4N7pgkSJIgVAkC6C16+cKO0VzJbxHZIcNF3KCObF1ToTpcHxiXjt
5d2wDDrCaVhNARmFvsVegBtuA/gxC4yaaosovwwwoewV0Q1QPPiRL/FVLLyM7Z3yJApokVfPP0mI
NSK6KIC+0wZ3D/LwIMZGAQe8bIokdUfyBPi+gA2Rvn3rpMA2LdxaReTcrjfBhfTxXBgUfKLtPPsu
7NWuOZFI357XNElCjAelaKGYhDWrjwIngyI/0+kiWAK2fDp8O60rw0GfVfzFxkUWYJTQdliv6ht8
cjnywTrWn7T8WukovX6F19zDKZ8PEZhIafSWJpzAaZsQ5hUt5mCcqp13eFastyxY92NSEBwV3JvB
L96ljbKZvTiFcNQzTXSaPuJXnyZ/e81toc9/yFlHR0WYjTXI6MjAL4572s0QPssUXH3ywT4UVLCH
PvqZEuI2onn+uCvD/neO17pPAeST57XgICdnL8b+Rx4ht57RwR9YNRGFrfkC2MLf0XxqO1T91IES
0PYKUvJRJaTSvwcwU5Zvd48FPLPtiDqf60M+uoE+XxFspKZzJwy5HGQZR921IKc7g2HcTZIZqgMu
F43KOAWxYtO/MavIpKGSdHAuVfCVJuoT3TwF0kWH0pBq7+9x/exdtDlMo+xPvYmotY4V6pBFSr96
o46AzuAJk0EP+mKBSnUUu5WQsd6oaIZ0tjfKwyz/nCFuuF86zjSmTwykN4M9sXnkqUx2m45a5ZFb
Pqou8rNAAfg7frt/VDusGjSvJkw9/LakHyftO9UBl5XzJJTFaI5OYPzVtr84BfllB2qsgF7SwLBK
gdpNg6Y76i7IVBg7HLUNgCfbenM2UmrkNLqnwqawOPhosjQZ4HakaeHFSDFld1maX9bRGIZkRnjI
Y6bur+yBIMix+eLhwBpjBBwGonDjB3+BwriWtjPCUz8n5aAwzMJLTz0LWXAvgVFy7kaSvjwyhpJV
NbC00SiX88Oi492OmnQ5mSjqTDc6YUyzR3ObtUwb25t67EfBFb2BxIST6UeTV0+ajGL6JWHbLHjh
yhM5Ky4GKvazBiL0JIq04VhbrzRdF3EQRQYuyaUzlx/JEeiL05YDwgCuTN+a8psHUhaZUrnCNyrX
eC35sLnXSWFEEx0QgJ7M1hN/cSRdp7n3yWv8yV+0GtmIs1tzqPZxx+S8GxMBHd60gDx1y3HUQqsW
Ij/Jsjp9tIvMfxfQ6Cc/7Drc9KxZYe6XubVc19Aqwh2EweKIRoS46wp5zlTSRVzcPJMjIAWhVOPo
CybdrJdFBlup3O+8XD5+KUXAfN0d9FGNfy7q3BOc65N2BPwjUuyB87yL82skRcvJ73rU0u+6XbPY
UthRW6LfR9h6geQEARLwPM/dXRdafPNKG3Ue2zyliQdMWsKLr+32lBMeyOBuq4PL0XptDkP0Hmhn
A7128/sN5Edi+MTAHpdOajijroP4mbuand2/QTGBzO4BEg0rj8/MIYXgOPPJDi6Evtgi/zTokHHv
jDs9GifJkVA/qRe2UeMaa0i1RsoaAudvhbAmKP9IseAwWo1yHt9Z41EL8CSsqz206AKvB7CBu06e
pGHQDYCKYeRvs+Y+56s2Oi9RD4cuGGNkodWQZud3L0a0wgax9B3DtP/awVXv7RMOpDREeYhZod1o
pI1ky8lGx1kRjXJmOM354i+FKyCePBuamf8uuM9B3cDj98oq6NUXNRxhKJlOiw3f0KRS1EuTa2lD
LgDOgMurmZhJPGIp/OHHIPflAhuyr9e/TuUCQOWkoPBQlkPlTRcW9C7KUjTDtzRhnmXi9I5jbXxO
8qrxc4O6sa2pT4EQm+EevCHIbCpJccNHm8SXCggoh4fB0MBtd+U/mP5E7MoSlzTgkvmzcSsMTnVQ
ZqrlsSidem/QQmUhj9PswnRbA6pM4kI8gVK/K3KYvbIuVhDhzZ4l1day5zRT+OZIC+62Jom3Hwwy
vqaoG2RGXdGhyAjbjMWjFH1+SGNjBFu7pwSvpXBDVpoEv5pGHKyUIZRHIfu9Lysl0LxkxXe6P/mo
tOey+ocH1MrEFUfCkJcbN9DCDOlMVO1P0DP/fk5dAQbU226nW7IQ9G3QuMFlmFemMWrBo3J8J3wF
CTPoDnfdqTMoaED9XICWp+PdF0cMf8aOpPC+X3+LFmwGRxR816hhxsQzD+YLPUo4CHReXk8nIQsi
IpGW015MtZhlx+xizfQwUvZd5wuXyqiE+bHeKuuJZ5y2/iDSdnak+7hE0Cub57gOzZxKB22zI/kK
otqKvoasGmH1yWWml+YhgiPISGSu+97zUmsyoK/BEuj0SzDYY3XBfqjxBQ3JevqRiiQuqjnGNgYi
UwhXDFmTjm7V7HsAB6tktR2tJ2yjuqqtmI93ksuMvLvCfGLD44r3ACSOA2pDco14J//QwXuPTw5s
uVC95no0jI517mE2ma82zOZ/pltuQMbTyR2q3bRS5gX7bKH5wzYLXigMIFCqwA/vbqBL/IgH7sUJ
IzliG+bks1N0BN/5ID1r8P9GPKgnLi/mg/uVbTgs80vpMYYMs9YYHi5nCP6egY0gc0FGf0bT5Hpz
QT68QKo77/vJrYliIzFviEQMZn35RP/8JcZ33vB3cMD/bcLcMxw/mvdMpQddaGqczoI9hI+Rb2uM
e9HsDm7CGYgo//kFGbPZ7UZhNuYCKrxLRIC9CZyomZ5gldXayP07CwSRV2XeSlu5Lkq+68m7WhiU
HF4JKFr1z2OwFK9C3Jpj5m7Jl8/Bmf/uNjPe8jqppKNYVDTSGT15/bpEJ+k9tdm1K94ByYlOw3qi
LZqo/YMDuJ5t4Ep1Ray5xI8SzPXPRzuQQv1e3rV1TCqv/KkV3tn+h9UyFdS0cNd+TpBRWf6zq7tm
95kbw+eLS+qr+chZQ48YAK6+IYkMk9063p2OCrQWgqaEqrTZRN6I/0zIWHVna/AquU/vkCX1m7Im
N9EMoFOcE50yDgqL3PkIxfZBN8MGibYjHhZyHL5qBWQm/nKlcvsgnCBrWBcvkRuQWFXGYWv+9mU7
BABKuUTf2hsa1fDfOiMYztieRkEFIKyO7qnsyggPr8T55WeP/8DjdWphXk+4G/L1OSG95skALJko
+WA5cOgZFj9y9ji7PHk2WtGnnwwdl78BDR3WZKAhCbxosHW6+oVxUejUm+Y9m9GdgiwHPjnhaI7j
+VuCE2PyZJx3M5nOfS+Q9N+IcM4UY1/d4n70Rkom4ou/n1UCSI9xfiNXBV320D5jByBvptLQ4SAB
c1QPgFGDxU+c4GmqthiMMq3MSvQBQgPWHB/UIMBxkEJ9e0M7CoO2LE0U6Z8XZJiGwlAJQ1cHmloN
9rwV3FQTODZvwJWo3pC6nrXd6OpZ6CFHSfALOXN85YNSwf4WGuMftSzuGXQuyO60hQL61mroqLba
6SpEjk/cusSIpjO9EguNKCMTnC/LpPfebK12793deH+el2J74QfXMGf+caTx7RfJVFKzHcs2kTds
eVR+uEAnwU+s8Lrmrb53X1Pk5eRm+zqVkw3ZZJNd8ky0pd9XTx5oMTDUMG7B4jTSHxHQSd7S2hU7
E68qmzPymVc6JOG4a9ieTMlH4+939sBqtk21Zxhu5FPNXO+UNjupsciS7Yy7C8TGW24KuS4nAMF/
hVGuuh6OjuGfLELi8qsx6ohXMvPy7AwauvdhudyXJcNa3Zf+sDeWS78DnzFbx1B5pDg5l7ua1zu9
hH5Jzvx8oZhb327gj5cVgrX3DIIfU9qR5HcWsW4kZzPfEz3eOd6VKazjdK59079Na/CtUbxJMUYS
+r7Kzxnhlvzvqvg0aWgdvKTDKs5ipkW9xClxZCXuMxJGTlE4qSRYEk8guODydP/bkV+YNvQap3/G
ooBr9o2HJzf93vfTsAiJTLB9AF8ATaJeHdY1E6cSfRHaiZtPRL87M3GyyjF2oZykKp8XSM+sjeBL
bIhHxb1y6P6iefwvR4+K31L9GnoMWUaEprYc5ItfROhDT3PJYrrJ+sCJLixAhu9BoTnRM7B4SNDt
/QNfeO8pY1QwYDCy2Bu2KPIw9KndC06Wrcmfs8JTc96VrKgOcehWvFGMoaBc5ZFoSftX7HTG3GVY
bAjHEFABGIlGMDBHfVqCoro1T/kpKsZ5tci65r4FhkFCKvqRRNirJZ3+Pq7sJzNhYOCQtxs9atQY
dSG/mK+D3AJQb4R7uI5GtgxN8eFI55fKXrqfLzAwp8xJaE4pV9wgk/AbUn3/0uput4YcrTLY1iqO
WsDrjDo2gi/rWonI0j4VeUdQUN2iy1oOZfzIxx3nUFUZcz+J/Vd+Q6nt2nUKcS4xytN5uIPlJzvn
s9mTwWk8eXMYEuTdbLyx+9ncXS3tRngoSfrfL3hbC7epP7IJoDsOlvKYUgaHQvZ08yasx4nsLxO7
QpWgmMTq5ZecTdNs8c2EJDa66JmYX4tj7zT3NqhNozx5oUH96ieHs9OPwEyDQXGluBgDsnXgRwL/
VwOZDZ1mhZdfWm7pQO04G3mWQwnmX/poRt1Udp9UhUqeZD+OMPGjnsZECfNRK0XL5OH9iybw7ZKM
jXh0+qD9x2jhSygNyJYtxNFvIsmF1ZktpohRNNBqbYaTVHudq8ztHF78KRbFwQ7OnLzCIj+p3usb
dBItQLUnFN4L0is52eAkxzokfMn4LLQ13sHLnsb4tTh+NbH0O4mDXbdUdCSi/J2RrR8xdQfcWnPq
FYnb637ImC0qocnImACPuONgQXFPyJ+i7tCXZ8wdZKNttbPhdoEDWb+raUnUMZS+7tcZJm95813O
sYW0KkcYMJVxCpCeI7k0Cy0bqh0ehS7by4OAEu2n2Nm6C8RCSzcVmb3TSHplYSUtrXxAg2/YTi4w
vk7RzlJnTssixEV14cbGZE2MbWh7klRKtPovDVPD+p2TWeqOmVHpQf9gweg0H6AEICHcmJaPbnHX
kVXAtbDA19aDWDPfYl31yJLyzIWj5WeDopU+aR/XxDnQeqD17SJM2ShQUyo9QyWqtO7XA6keM8Qe
8nB0ZZ5YSKAwaK4La6XVL5t5D3e70FQXpAGzovIs9OkY8vPog9Zv82qtT3ImDU3MvE8/TZOP7E1N
p5Ct2E1LoKgqkNc45S3ItzeAp54GXzoVEHU36BeMgB1xJuuNPresvwJRUpYtFCnYxrlIwvhuJzbA
Myg5+y0pnSg/+4g5lYKG+4aGBa+2EPxrBWtGLhYbmVon4qXZTdnEibREmTKHHDE230iO+6V3qCnp
tifMjyE4Ncrw8kn7mSw5glGc28eExNk4fEXvaUqkjz4leOEfhWiMYVTGb4ysii9SyNl3y+S6Lbrk
GLez2ectyZIuF48Fqh9WsUZL/ogTurXtmOn8Q9Izqj3/Woc3Ydnp8CAuXfFxovNjf7PakIvTyI0n
PVawzsG65jWVcrsA3S6WQP+Wndol59cG+WTQj8GYCDDjpMyqAu4blSdDTBopelry3mMVjh9RrpZ7
74nDtbIjW6jvhZt8zLWXFcm+4A/vi2Er5uN2AnnSY8ciqucg+IKqJ6qICGROPqCElYM34HNO06Tg
ceKIyaz5JwRwnlcDomN6CWWGIJH2ejYHHnG03kOoN0v/AwVz9BRi/U5fBdzBS+TbR5X97/Jg+V/N
NAfl0k0yCT8yC4mN2K7W9ESFL0jjXP7zC0g7vLJjn3u3qZ4pC7PA6RGU1YaYiN5JpizCBSEJdI0K
zmhbJZJk1G+oaQAgjJSHADFzvA2+G+tbVOBLp3RL6pVcmr1Z/TRosBx0I27+7v4YgcsnUFteYmnj
5i8ao61f6WHdoEwj3O0gUaFKFb9J1e+6yW5Kmi7yJsGYwytXy7DkBtQLUCuGNjLCcQrSLBKSAVhT
QRpEp/h8oDAd1HRQFWHnvr+vSx7/KzV84SMGbuAeR6Hn2KcfdarIoud87VKXHc/+/cb67M2HJZui
1bgye5OzmgOUZX8A62yo9iJ4mBsLE3MN4rUJyNzjFlzjSwXB/iDEjN5VWcAop5JYSyVq9zCRTfSq
tSE/FJ7QD+7EQvZ3H/Nvib808W0t14KO7xRB/8koKLtfKqF0LxkL8SBL0P82J9gm4o0m41LngWaI
u7WcKZEDURNCpv5YYTuZG7OCsEE2TMri4byaPIDHvfJvyg3fEGYduq01y0zLqC81+X2cg0PVpEZN
ntnQjsrNlcJFXVl8d0IA8GqMe5xrwvCsR4arIRt/6/2FU99AQomCs1nYv9K5o4n/Q4UQvjCxSr5D
GuMRETvmK+Sw9Cn3JqTDwOQrCuv2Dx45bKqi4h2QRTaZfb2LN3RQbuTGY0gD5y5YKfI/YJeuAaAt
wQ6GK6YAhtQt9n3FSCcvtnokYlMim3nA29RgFtYYx+Hz3pvA0yyIM5YwvdTvDmoOtKR20OmSKTZT
dJkGE5AGQiFkSFSyqnNHUNAAPhh7zt1RL9LIHnDYg/HXCvzDwYmUk5AQ71qO0RteQkkDybAn11FY
vw0RC+b3MDN2jOHkxrF0zS9/TlY/j6VrB5tmgJUmr0KQwDtDfHMO3yOxZO5I+SSWsd3agYxP97yl
nJXcs6LbJH+cjBR2Gh2B2VD+Ul6A6mckS/wbKxxXxjpoT31IG968eJo83VZQpIJJAqe3VUEVUXHf
lR/oHUfewCeJ6HIbxPZ/z+bcwAbpQDriNhzfLWqdByKo+aw8TeebVGmw9vetwtFOT4MFobgxF58D
VtrVEF5m+yBSYSEJgIugcEhGu5oKuuZKVV+A7P0G1XYZj4bi8IoW8QyTBwKP/qHYIStx+UIslmU4
JIDgzJar0p90/SfCzB8+cNHNhEBCZFChE3AgljVapZm3o9nxv7ru0tnNnmK8E12gKPhKjNzyv3CH
BBIUXbVLYOfnR/J6V3/l73Eo9ycbyqsPbfv90IJkFbJLkqxo+4B8G5yMFt6KbEmfgk0JuOkThrGf
slvCTPq3vUP02VXCEudk986oQdQqf4nI5UTvXpKdTxOsr4c1gW6B6hsO+vNojuaf0wIchOSpwGfC
4YLzro3PZVQTA9ZU/YOfvTksW+T5cdhCfTaC3r9eXypohjQYt3fLP9MbEJQ+XF2E9A/OugyPplgK
xjMdoyzHKvNHWDPA5Xf2tG9pV9PVpZYybmsOG6I4LsZloba3ZzJaP8R5mMdiU4omxCUE4gu+wdPX
s8ob0TbuB6YLufCHe9Godyut7kOUrMOSiRVYaHZhyPN64i24ker6T9Xj9WN7URJ+OVXfN6GLW7BM
VyI8tNYNUrZGzXTaNQ3t2O09EYxOn9g/MHN0EWDMBYlib8wNIixYUNDe5j1we1TWQGlWDtQDIor3
ipxuaFVrMAwG//b09BE+0Ehkm0I2mrYmHHIbk3iL17H+9uBKU4Uz93M7uxnmdPoLksseOi8x89WJ
8Opctz3W4WO+A+5rrjwxDc0IrRx4GFagc7urQWkU2JekBvsYXqcA0APO8rEO4sb52gniFDrFgNdE
Qihoex9e0qnq5L+GjSaD1OFumdyjQR1MXFXE29Kj0b3Nbp5O8FMA6JU7Zx4UYqRbHQi10KNLEiPq
3EpgcUDSBOpvuH2/XnJkuBIGNh1DxqTCH5le+VRr7P9+TS/X1JV+5KroVNvXwyOL8aDVD1n4+zB3
HGI7rub4Z3NsvqP8hScEqyrgZA6KlG5DkVbw4ymZyHxO7DAl+zem8Xx6mk/O7gBJ629905174Amm
z4/M5TbsiJgdaHQJlnqe61veftD5Qj8l5X6IM3lXQxajiw5C6u0VQ6IKcUSjUV7mjrcSysz2gVcy
WVg1rBWwXT8oUGtP7ZNekS0ps+iQIcKkMMEeU4MXYldr3cwlhi09jCvRTdrYi2xuiCtL9PG/qkD+
Q5mOwiK9iVSBIhUI7Jkzzq8gpupzEI+DuXJi/jVfsZq9hslgQaaKjxZqX69HGYFhMMWQqWK7ec7n
Oey4XkO0P4ceRcjeMw2t97ChOpaYys/PCaH600PiRanKsMAv4Q7t2qF9IXK9Q1o2t0LF1p02lPy0
5/bUzhkUypXKNIy9o3sQq+h8sbFvU9aLZrd+wwkrlJPHi15eqQ67fto9a6+P/+poTtN67io+rhxl
0d2w3EAia+pZXLXT5MgeMTi3/veOavkeN47yKAl+opwbi0IrR4qNeNGejkELkaohGV1mXzyTNEMn
XOHg4AVneiQw7dWPgINNZRXR7TNVvZs8l/rK5Zt/ezNwvx759UBmjm30z2KJ3/Oq00zZEwzsFhwV
HDC+yoPhMSqJVGYmhErs77cuPjd/X5T3URMRA18nCB9rFKtymGQ0ioWj/d45rYR0g+AB8xkE+22q
i8h41jNyEJ8mxrfcUxlle5z22nGKetfS/sfB4ByNMAxbRsWM2wUp8uBtMzFoUJScCBOtm8yFxVf9
i853Y3dkWUBCrsD+pTGDP7qmefb98mqpewjxGWfjRLb+SkFO0u6cNby14Dzi2/1xYYk46woWc/85
6RQA+3DQIEkx3RjaBtWVycrGFc44sGEcArP8Oml6WSJaxbKgHJyEFtL8Vqd8JNiXwEHyRKFruzYF
BXvcPJxNzlQujGCJBoudt9UnxUUSZEQoJ1oJRg/FOL+fDjpQKsZkbGPhoSaf7YAjvV3nEUBiwWa9
F7BODmDl69CsdE03Stks6TwwIPEshhiETjfv3aVOgboN4+FJeZOxvnhhRTfdC0tQrb1U4o7sOcKy
WVfiN1NkLrthjoZYMnQVeEMQeJT2zBRaj24bz2jnau+zNZAcXdi1/Pa6bXPMbjvK/8O+50bPzZg9
Z/uiYRHicqqVzUzdi+RQnJVktWIrTUm5iQV0F8i+8VPg9zqgHsl6ioFohTrNbHT/hsjefCeUn7mO
I5fMeDCboJJWu60NJUZBCNJs55CK/rzaANeDWi3ZDML/YISETrb3GKFD3/9gudxtrX0+++X3bkfH
ka/9/5ob+Hf59IJV1B6SBurMpJzyqWTTTVf3MXWTUb/Rm9f3Ft5D9msRcZoiKwny1DuhOOopeQLm
nYw4ey6bfPG1PnVjkb5IWrzB1+zXt7qR3bl0C707+OEGEXP6rNdGqcwotlrL3aseg6lbG8flucOE
xIlg50cCmsa0aRjiGs5vHprIdSrkY/VUqG64xlHjtHqD0c/qT2GWghmgS57bcXdtR/wWhSP7Pp7R
I17xQSYYPFacEKrKGslNDqNNBJdYyDpNPHiEXAVeWxS28z4NT0e1v0QgwTw6nsKP5lHI9Pfu6eOO
m9WMG72wXBR8vx4tEmmQjG5PlL6DOWwqd7jffi/dlcE9E991nZfoQh6e2p0y+9uMxl267otSoV6m
TmfY8Z9+XYEWCHWuTUH+DWUTEJ3dOW/maw+BgLGYydF8zNjQeBytZ5rpFUseM/bYj0t0593dNGBI
VQa/0rZrUsVj8Kt+eEkCHkfZdoBlbnmtvdJd5Udof85yqbtX+qKQz5B2NTYeGmZgv/4CpmgSfjKZ
K66R4vvPEQH4mSVF6+oCg9uZ5UGl3ADbilR/ixWCHLjLRULrP+7lLJbOoZFxjxjBu/4sAeFsxW4f
TS1Vy8UpeplOhdXpHrIOCS2DGMEchFXf2Lkwk7PHS4mDPwvfdyIqOkE0KeRO4Gw4r7bUbIVtF2AO
/LTowLV91twvdurHxlBZMyxKO5XyXVtX4F8D+MW1f8gOey2XPYvDB+jAMOzVGVM4B/ObKsWeQbXP
Wr0q2dc9fbBsdHmU3mu/EGO8ze39/H24/WghcwnMIQNswIeclcpTuaRoM+55lxHg/GHTWqSd6q/B
kwieur5CeXmCx4Gayi0ojt/FtgzRzMg8KC9PR7N4z+tK+82cS+7DcvQPI/3GSQzsfY7Nhz6yZcjY
bQ/RHWjlF1xgavgcD+fwMSaJgS8MWENbFCc8u/Oo7eTIQ5W1Tl1W8jCCgQTaIhqpTXXMkOGCqOuV
i5irOOZ/SGqOPHT7t8guQ9MspzhX5xvtsTrrugK/qo531qeqhI27pSLl6e5UrcafJEeIT7pRrBe4
PgoFAgqEYENEPf+aDsRtTAKybji4vcCXVthBShNdeVcOnajOPbzmLx3rYMrnFSGov83HxMKuzc9U
I8lapZM9Mhn7KSNImxRpjXV03YP2lpBCO3I5Fv6d0rUtUNYC/PSMgtQgQM7gql4uO/rr8T3PcOxW
4GZzaYjk11zbkbKUHQppMhQ9FwHicGVNla78V1YmRERjTzOB1ocgZgS2bieOY3jd8Fgd4j12PC3Z
/fNZ+yQ/FryGk+gWOAa5HHRfHCwwDbBhZJQOo9OqGTRu2Nvu/RRhL9XgE+8PYWDNkL8REDRvygfk
3TRUoPArAOLAkaYnWYgNErtB7lpgYncGxU09+WpYBc5VVuLkCx1sKrA6MWhk8gUkcueqTyP35qux
xOXMqcRSdmcEM2NQvT7SvrLhhXNsrz1aQPicLL+UMqplPKYiCgmGjyPQaZR6wZn2zs0MR68bB/tN
R3mtK0j3km/k6vUUYhMstO/yzno34rfTyzK3+9fB+glW1p31A8F6zC6EijLZPIIqmg2f0f6vGZVC
UOkoAYOFUwCI22iiTRLX+FZ1UnUVvEmZ7S7KjRu36/q+KrXmseFbSqIPGccJEBtF90ic7sLnIEUG
Chk6FDUliadtvwuijda3V2KeKglzCxQOB2a4SISgoYQieApL+8cAGZl3RpnvkIoCZJSeO9r4kJr7
EC62LNqMUcm2xHvjDULE+/0TILkBNfuzARhgUayQ1+1BqEpHGWQTpWMXKK0+SlTlBVb6vd9eR++q
rhNQF/KkVla0evWWg58RYqS2HzB2c1inkVTeJcIxpSYKmJf8khSsuDY7JXZRx8m5AsVR058qLLzh
tDcXo2Sg0YUpoqwfLmMtmfoxQsMf7NZ92V3KIJqhit8iY4JuKhqvW1wihQMt0kkL3+gyJIRW/4m9
chupF64LMbbDVGARduBRd3OXvZCZ+/wyi0NjN8mmPnIFsSnpj6lFwHLI6gyTimvMOm+7vcAy95nP
V9101qYvRWRkGcHDCOmGIMMSBAS626z8jOWuwPitTchBEuhsRhnJQHcyanMFBU1XnXUqSmaOs7Hh
SVD5O7AsxFr5OVgBjQE22P/pjI33Hou1ucz5tWbTzZTydlQfn75mSNwvK0DPUIeOSbXAziTliI9H
HlP4Wdu2e0MhYnlTm/e2jXJtFIXqaSijZ2EnuzV9A5jlZOKih2u2aK0DNSS03Z2PzV/D1Ovpw7c7
uIAi8GZcpKxAyKpJJC1SUiBr46VPoVeZwHrniuFdFytxLe1pRMNAv3W8ge1hLXsV5ixHH52Rg0QH
tzCNmyRm2GmutUA+s92FR1L7XMc4b884qHZ/HXuQ2SYNrntYa8R6wajbfizhSKXYcpifXUuComh5
6g+eaFrQrMhn/uEd9kaw06qlhKKfmD2pC2+5ePcjnFBbib41u6ryFK3q7WujFwhG7SlNUKRcxQXM
HtUv+BFdlS0GPDdNzffFY0Zyi/CzN2BG5M5Fe3Ghe1CGSIyFbxdXsaAa69js8QR10jSoVxKZhuQt
of8OmVwohe7f+d85ZF2mCjyOxeDowA1qrGWWBdazLn0Hc5M2oW27d5vYpZXuCtf+KXUsAobl6T17
e+B2/tLkdso0ElWio4f0BpLjUxF2lk/gba1dx4oB5XbqMoq10CIxnEp0gWzGL22U2l2Hn4IaFatM
KLvNnGva2mVrpBRzj5K6WZiXycjpYm96k2hO5Cr3RBTftEFKcZ9g1q2NntAbWu+71UeWcjXk8G9c
e/HbzCHYJJIhBOmT9vaRo7IEGHLBMyo71pJA6HL2TmAu/NOdavCIlg2qrDirAtHnVBnU+OkTo+lp
EJaneuMJOTsqlOl6yIKS3rzypykFA2XZD/GRZsjBCgCKWkPW54z5X/ytTMhaUWs/wvfRz18nGaE2
7RYHNVHSmN4hnecL/5HY1ESMd2uupMGO7le6uK4Xg9l3HbZLVazCikICjCuTFC2Fxfqnm9yoxYqb
xEIpQ4P7knn+rz/xUTS1qB7mis6LAVtczLDix6aVsk+w42w0scy9BCJn7r2ttzK9s4rJzp+5TXKM
GYEH87IPKSe7hXfqfPYO7frK/fiYh7qhUsSCQcm3olNCVL5o3yZ0kEY1d0Hu8EWAGyENxTIT+BXI
bWzrfhRy2EVq7DvbNzVbLmtf+zi6cavRaZnfAStS0on42iU7yuOlbEhwPz7R4iSsFEeAM/TvJkI+
kmsBEzR4URxVagSXcowggBqiixzIUA/3qJ1nkq7f2pKjDwhIbayR+gU6E4+n2+GW5N45hjHa2Rq1
w0KCap+ji2JykdRuRAxz4eT1l8CazTmOUvRKCHg1uiZ90w+Etzk3R9oOVx2SciXPWpG+7uYmMYt/
DhAeYZJCm92ZJedNrZTwn4NMaUF20MIYLSVg5rlPc0glfSn4MAK0AtbVRXdv5BXWMwPXa6WeJBfC
sedbvGZknxoJjyxMmzYtUTqPOD+zY0RvjSXJBDaCy99Sfo0eYKnD4cEvPg99PgVstF9AmXAXr5cO
G+7u2M38HWkpjHveXGzzDmQGOPIQwHzD33/eKINQLitu8qnEnfcxYBvQ1x906d3R2+NaZMOEX85y
7BohLnuSoocygUAtLHwa4t/zCC3T22rSnKlVwu+uygSG9aINfFx1HkejCVM+nyWMD+CXq/uAkAMs
cTQK0uskilECs0qHM+PW3vkTEJE/vtEgzq4vOTzuSFKxPd/3ZneMk/Wx3rQWlhSBKSNC2QwDMAHC
rg0IY5kaVqFMUe6AtFGPypVdVdwJJK0kv+DzB2CnA5ah3W03rCQr45VpGBd17T39JDQ23LaJfGEJ
L0pb+m9W4SbvEA2i6DzVg3ah2/Dtar4L+DUlOIqPj3SKliPTAlekcCRlxM+Q+TJOydEYBVIo+hsV
Rlz7IXnxBuV18l6M8NjSYjSic0EmG8tnwcTJFKFp/86f3d1ti7JdgLUVR5KPf115YI8XyCxvpZNd
KEwyCe9uPOygfqQvxAcxDSzcjmtVcpOwZ5gEwXIbl0HFdmW52uIIXFFqB55lzs5jsZmMBaMPEnkt
kJI2Mis59eaGaCev3Z14Zfy+ZPm9WwybAWMbCBpuwqUThGMsDSstm/zTxly5ko76NeReYiobJzaA
IAdUsCWlQtOnht49mfYmsqcOdB7Ime2dshnzzMbnTf2dSTdEUbvLdiD65+lT06z3sVhKCWyJFO79
Vx52s6fVvrq1CZpx6dfWC5EEKPoIQJFdm/F6+NrVi8DHpye4IjnOk6ECvnXWCFegVdEA20X/kfLK
ECbr/de3eNFvLbUd4j3LnXCnd/fXA5JymU2wJySX11BEViuO3CoCMDXUE94aNNBWrq8DFQ7tXipm
UlpRLLxVBH0CaKRH2ZHiHOyJ7seQ32blzytglFkp/NXYQC5yAOJAV4mCj5UGco7yqSIk1sstS5Fz
0f1cGjWDRGHYEkkLBam7Y+VnGxXRWFa2ohDNALtJRSSDhb+o+1PicOVpYS76uq8gVoDESie9QnJq
sxpma/D8aMQBCu1kxAi4x1sN9hvT2wlD37VUpGnIHHj+w0AzcWO4RLhTIpm7FcIZH4qsl6Za3QWT
q0ZjFRZF+rmb2Z2fF2tWsNhSNrUmFH1dtnaEHf8h0fFeZ0oo4FGoZIrwwFPiQ6ifMtBHBWT+4MG/
T5dHxdPdrBRP+u8c1RJ/KcdK7ayIT4+JHbTR5Fj+YB/SpwfLBfAbigH5j5s+cjw/r2ycmYPxv8oi
zyvLJ3FRAQ10YkTRpcjhUYQmtJ8+HCX1ZDCFnZG0VYR7+PPST/H67KCjDL60TGD26rRbY2Mzm3lw
D2+8OZnJbIKVz0ctDh634jpfVKTB+5kS/1R1bF+puaRatVQrlq1XoAEDKhq3TJ+eO6XNnTwqLRaI
+xAG9mgdf6/KbghWTLjdFeijCubYZGB/TMfJiTQKGZr+w2GDDmLwqOwrEi8xkmEqNEBOovys2XjJ
pmBur2Uhu3V6Oz9NnrkX8hZKxxMbkb9WNrCJyO26DAGf6UZ/wyWrWDI5V2Y7kb5jLBR/4gJqb4Ll
A4JVAamLfCWFjyOO4C7hTpv34s/r9wjIHHfrLMers6MewmpWU0FvffUJw5jGIVvggB+cmsmX5LJb
99HeVQSK8hKKul/JkDyZdR0mRQKRNDmvZoLxelyquojhhQQv0D22KylcHVLvbi4nwJMxXwFV+SDB
SserDClqmEH6So+edK6L1H3a3eI1W2ImkurbO4TlUMxkrbmBItONUxJ1WjPATKhHX8YSsSJGIeCM
qXPColI4HXf1Nb+AClF//owC3SPvYWlsJuhYagAHIPDihC+gMYcNcjIyeYzJ3f24W/FPguvCPbxj
664HEiXSPJa5WnJE8WXEg6dncYGMZMO84jaapcu+RkdUrLKAvNViwPzS6qSs6f/ycon/byY1vuHg
hYc1HaqSO1mSpC9IVY5nrwbl9JVRQjPbHOKOgyzA6wJVBxOO9Y7HnDVNwkgLIPtyFWVMQrZK39MZ
RTTv/nc+iABNeV9bD8kr+ThMwiKkDbb2kSC/zwT32650g8xf5jEi/QOjl0M09rw0dSCcRLpH811w
LvTyB/c3+59M/HSoA4nrpJVHdknyJfmibStVpmm3+rwdfxraTwAi2yW8EaMXNbHXeYia+Rg9q82i
zGHBo7pQGgn+Zl/uWYYqCNYbhhefk0irrCSo8A4l25gfnKzoLiXpRqK6jhs+SCTTHXV+idNcXyoZ
Qe4DJC271FBBZckuMtJbQ8Uzpm+AvQzXh8k09TuH135DHXOKa0lyGLxYEY0ax5TWkgBdzxKvGeCh
iEpp6BvbtpAcfjcjsI09K2cn2yh/KJ9umY8euVHxIYbT9Jc4iehmM/Rt2bHlJ4jv/bTN88VB3wsw
4KDnMZeUNe1i4XUbkTWUa768RkxgaoCJy4hRdhou2Heio807q0xpwNOQjL0KT1DWVB34eTDU7lch
r+Et8VOWIUxzFuvIf/7iPme9QxEvYadj4K2IGjFRNOK6X17JeMTRhZBof8hA/HPBXct92Oy6WEX/
EbcrwH+HHjueQSFht0ioKaL9yIaXZMVi1EUn/YP/S4yUHeXly/nISbhVp1JbZ0By8AQHPTVZqUDL
yl18hAHNz7OLZ0T96hZkWYgpAk/PSEQS9N0X+bi7wLKmTrie1JECi8ahImprBSfsjuk/q5wRrSUQ
o37fqvWUr16nysVkCVITYmrWj7FDmv0CY2bP7mtjqR/OQFtrkZluy5wHg6I+/tO4UuPd6sWoG3dy
b0gmmIjqPetEyQ7nzI9opswGCO25gK74JsUAud17KfVChRmwz+nln+Oz6QWhqICjN7NXVAzqBP6x
JrnFZm+PAvhHhEUNfO51+zg/kbsg8atg/S0i1xinbtiQNcxPm0VK4IPAgAdkHRkQuxaoSUv+ok8X
04TsvLQ70LwEgtYAMOF2kmp9F70LlLKBIBtJ6ZViDKrKK+qJyK5iNB+fgaFXfUhumTZDAPTQAV4R
eQV+ZvotuNZS7cN3ovkQjhfb/csfMvMXdlWIx8lYJUB8icpfHTVVzhsu9BwVszfydUAvXnuVccFt
bzyHVRlTjyA53MAA/Fgv+ZnW0mMeJ/fk5meIHsFTUoTltzSUpI/1Q2N1Fm7f3cgsUDAraOwB3n1M
2miUuZqXFPED36cZQXqccR6W86uou0ebyusykd0Cks5QqDW7yzREff27uCr3qjK5bmeWSLdBe96O
D3T7L35xQjMB+i6g9xDcXm3/V1aNUJpgaQxsnN6w3GOYxOpIshobBXt3yAzNRqNl8ByAdtHIW2ux
tz+3OKDLapzGSVUNUO5uyvRopDsECUJT7L9dsi5jlPsuwWRZOSgmnRQXbpUJvDdVaITDZ8iBCJdF
sVTktqVCDOiCtqP9axiMZVVwJKp7PE3kPtTIgNjlmJwLWYgsZBxBGQV0yb5mVDIrS8P/417YtGkJ
ex86xLpWIU1NnFWlNW1kUsxpnDlB4OWiIPZFS8VKrsK0wc9wbZC6uSWolCU9zxBGu62LcHf9TTsb
+m9XbSZm9Koi5IuztXaAJM1tQ+qt/aE/QKVEmSBB22kbDoiqyQo5aY7BMBfLaLrcfETRbrw3XyqS
P4RgqQTr1cYesoDgvAygX0I0Q0e/HfhgroK+JRW0aP94PBjYQ9X/7o9HkYVDiWqTVAnhGeA34KEZ
0as5tLDN/L6GxFZmzIIxe59SCT/PHfZk+GjafdspbO9T+ZfzASMG4Cyg2zbPaY9gtCdfsMXkfpu+
ecxY3aBQpXEnyeer6zmPCZH3xa2KVuciENCZNfDSldUlPqW6e2sTqgPKTLReGTXQBBQKFmCRm953
hglUbuYblla95gZl2ccr/uAKPrK82A2GaHiTXQNRe8coUlJhX/XoTTzx/fTs0Hw5v9JVH69+HsX2
D1vsBhDgw439sLA4mujHMKrPEWlaE/YfzENozC8XbvTcIPfOmpTJRqyufFPwOndqBACrTznLE5uC
z3CM3fRXTZjc5/7bVIQ0dmmCXUWQ7O3Jl/5ZKzTZeuu3JLre4XLPFDYpvCh/2Ai7jys26RonHhiX
38N7Ol4PHR8ES/YOuPjoTbbhxOqnFpdIvPsMUd35XIsRE4tLxa/yg4NNi4mFlP4nJ6ZCCG4QhQhJ
OWxcVQMRHkTH8CfkO3q6iLhDWS4tBjCbukU1Isq5cwxiEV9q3gm9D1iL3iFPfztNynJUgpXrm1b3
v18oUBe7Kv79G/T1luriI0J2ow1MQu+gFRmjX/9sLDlYwwsXU8imdaQMAiXdWVVmDu0w/Bk92sSs
JWyVVjfsOG6iBubyoWpXLqPcDycu5PqlO/Q6ibeC+zdZKgVXX5gHBf1RAt2nju9MNIFzly8TBZ/O
y9vPplWNdhkc8zKLtJD/cG30OfZQ+eiYzB9lexUQ90555R5CdXuzQvRxd8JZHRRt47jUHGM+JoaY
Aw1CH8njq+3meemkvO8f9W5c5Vso/XykWFQJp1AseDg/yacDJ70/brvG8WRJ3L5qUnHMCX63wUyE
qX3yezCEN2BFRn9I4IJ+YaeELi2cfP3e8fvJyyOm1HA6dTOGv1hLNg3uWw0pqRhso4f3rubW8CWV
ioiXM3rpaEjFZsn0n7Q1A0ze2mhk6n08rHfZcMwFvai+Gxcm5N+7Hu7bsOaY/GUOLXDD2hNTgDX4
rgD96LQVvs8nM2jxXQQfTPp8NTKn09sVcN08H9jAC+vLzugBs9ZT3bSooPMhcRSZkvz/W/CyQWyV
PgDCmbLGPrbKfRC5Rok5vWx/fEgqAbZ+ZfW+o5Ic7LOfjLjt9j5TNyeKiEGjUUi2/7jpZlNu91Yy
Y2Bl8cbWqDhrTVVUq41yZWp+EXJ23LER6FyKjbWHZiiUihHu6+XC+EqesedmRDj4wivqohIydvv8
Zm8yH+ObtaaOrm5EMTKve8nqEFl11Ei4ure2iLJX4NJSG1G1RaI11/hrJRnB8tklsqJAvQnGrkvx
owR5INrrmwUDrNhy2CZJAWWzRO2Hewei2LnLf1UCSb8xzFn14TE9+f+Aicixjm8Vjo4wVGi/X3lf
+BZIAfjG4iK6TCT0Dy5SE2kAyusGPfKpiG4kRLQFUlHc3LVBHBpF2IRYJkpTew981TcMuptLPvuG
j9Qj3FiKnR5EntxWv4PfjsX8J3aaaxnrvgYNB0reaZj+Od1v2vOSBtDAXfdvogkJjm2eNNKimVAW
xzSRvc0g9jivov/v0lGaoNCZm5NmHVPhxIUUbJWjHTBpSWq6BLbHG56SJ88iU0AYTJ6MZJ2Xj/RN
uUjAVTEvkj9uHO8YC1PUf+tGSGuiftGxK16JNBX0nlcgnaUJwP3LEf6qdB6TYYopM0SXu0P7WD78
k0U3qnb9T3Kl2u6/F6YineCPvyLSj5hGrE9M8aPbvHLr+QC8+fF/6+ZpQVnJd9jLDuOsCIKeoZwZ
rdV6go1R/ysv1z5+UKFcoyuyQdlSgsQnDC98jDvC2juLiCDvyLKE1wzqz38yaPZYaSFCEEeNn/Of
0vL7jrgq2JwVknq9WV/LyMYIsXUmNpBFWY2xU7uudfnNyGVuo1qDUpfbNDV3WZemTyuXWNyhPdiM
eYOYO2RRG4TGvKLsf02QfOon5FCm1W4E3zWOr45ovF4U7WfLboaBqG7B/cxhQVe50V7+aUzT9lo/
oyT9JGtgukJbwC5Mjv8gpMTdNxpntUEXEjXDYbuYNfXo9jvGXln9RmnOUPjnXpOW1Y0KsMc+AYUI
nk7YFlXMHxuUSGT+HRY6JDM+9ndwSMqkL1HvsaFuUR7MoZP2grUdK/PpZ5owX78gwTzYRAP9CGje
BeX8jGOGGTfztloJ59i8k0uNMYyPqiwNRFMlqxnh744VH/p4l3EIdHeBcgJaB0AUQntBhWkwlzBh
P7sdMl0D3miiI8Vy7QK3FwYYPC/R4MqrcapvHgqjEKg9qPWkT77rrLC+eUdpx5QxZ6M7LR2usn+r
6V+6OiHUxXXdoZkmUpIGMv5QbxTAgv8rJd5XguqnROQzJzBL3ToqgYVjXPymgABFpkFBPecaOgBo
Vn+2klJ8wH8mI5Q+QKChaOx9O6zARplYT7HavH8ldFdxeTjBYajSjdwyFtPslJbuFLOU5pL5z8l3
kHBKRbrSqWnMxKXWRuzVCVu6XJHuznd5x3bZZLGiR3E8MwrnsTklE6T8B2s+DiJgR6xWTSpcjjlK
cFVn0fo93mza9PHAqkzdNPCBu55dlPFgLPKKN7o5LMd9FWc+XEXRXGXKL9fK607kgNa12vVPen7I
XddQ2cwHkwswHeHmlZyc/DKqfWqzYm4Ui/mHXhVLE+6OT2VWE59KdzIJ0ci5bh54G+J5vmXmRsoI
Y+paXOWDc0qU4G6030H1LZOQH7ZIFSpyyr3esS/Cja3Z/PfSfxSlhD5EPFT1xD8WK7TCixJrTnM6
RxeWmCauL1pnAX4r76JLji135t3EbPXuPNaOI4WkgyG7da4E4JNVmFKeh5eiKvsWg8B0+Fk9C74v
12e+v4mCe7TkL0kCvpGdjrwisXm13RlsM7kX9NNy/q+lJ+GadFxMnj10AQpTcN8o+f+lqGgLofof
kNgm7+KAVh7/TGZB0KfhGqSl1kSoh5ga44wp3LF0y0EH54Pj8Lz67ShY6i6vOoXRXms3LCvVB1hy
Z3ztxLo/NCiZ98KW32Z49LiD009YgcZLRozdTLxSqp/GEoFCHySzrAslGk/ENRDAhpe8KSL7BNRK
4b28z4/Yi4jyMHpC/J/8tlz5lsz3/Tm7fWLptq5c/FVBmnBccQ2lszehrB2Cl0tf4U8BlrO5Ze5N
6MJpEYEQtOQk4DVdVr4UK4byKFmsFKUfLIM992RbNZQjMu87BkpLqwmjT4l/bAfGG/wU0QNDPUan
velygrL7nCpQti1BbR3sKHuOBbsoZ69I97Pyr/NbdTnZCDpQtAaO5HE1mhTvlxEbMrhf1Etdk+EH
PWrZovSgAXb6XWDIfzQxU4emaC58o4JeaGpynQMeuYjEaJjSAoqMbTjBJGRJmfgWaib6+425UlLx
e5DpRiziJLKH4Yu649gPLIfIF5vQG1rGzsnuI/w4AyeWK3+TSyEKklgjsc5xr3enRV8jxQpMF4Oz
c03oLhq37CVtKRMYe/9Jf3tFSq/IthD4yp5Kgbc2T89j3YZ7kOWI8D43wwmlTQe70zxqu8JFX24f
vqQbdflVtyKIyMBoiAzUnXbb0/cD7O7c8s5RjqHthRFWjKEJ9jFY/wESqwtqfDVF03cbMQZbqmL8
EyrBqaglJoAvNnM/cEGLEgCS4HL3nLGS31omxO6lnPnp5Osg4kn7uThmU5qDg/Vw+fSRQR/3UMHl
NftiYJGVSs91bWx+z40fh+7cQ2gbCO0BJ/HjJM5L6urVAOdpO1FKmUOlnrmDoqSKfjsDniOnzh6I
xsKtLdXXLKatb3ndPfJJvgQYGa96qcIHJDlgY7/wjFtzJUDFWhjTaMzd0SWSg29266mxhuEjWQg1
Eg1O7ySBTkDNXFqOG7R03iRyjP65zd8Ur11eKPlgZERTE5rMEVuJcxMWMggry3UJZWqGB2Q3lYlC
h7fb7p5nBioDqRbY1iklZpa1XQeZeIUW8e6I89f9sbTEcu1gWaCybWE2IC3QrjxgAGB4ZlTqawKE
cBhrO5rOQfHQypr1SPuHDlgXguDXm+fZwWMkRzaR8hPdrYYK0PS+dJ2OMUrxIVvXJhEmByx4CRcW
T+QujW/WjJgcItXY/FO/yL3EcEjNVm5pQrNiBlizYoyAIvpcJQl8mRiLLs/r2Ga8I72u3MhjwKSv
y2XG6jwPpDsD1TnIqnu9GkE3GgGNv0V/j7iZqmyE8fz89lpZVJ6NxklicYWeDtmFDG3xD8Ng8Upu
s10gUREbkIdVQ4M6csAAiu68kuab61L7nd+0CGmzH9Tkr11izX+xnaQpMO83KZoqUYHLr7Qt7FL4
P1Ja3xhTFcDX3eKzxWI+oxhfDeDWqI4qBi6B+T1xqe6RXioAGk5OkSFQQT2uNE7kfIzdlK+T5wra
78k817TYq3BEUHkjvMHSmD5TKehfcVMbpY+1HIafhuFH06vtchgMMkQU//JPjKu3p44CATZI3sbX
pd+8gEj0pUtusIMhKR4plFG9JG6m7ENrhBTSiuKBekNPlUCvmDGxU5QkQBKPIJsD2dDbTG2m2KvW
G1dtymbfMtfF2+J/tw78UO/QZC8hviJHp+csMQrJPLXznb7P5gcC71Rj1d1y6R2v5qzsVmD1u4D5
AQVo82iR/Frua1sVEH/e7PnNNCSMYcBDePXy2aSzbhuNHbxncG5EZoWhK4ed88zTnG2YtEa5/Pg4
0tc60w6rn91On9D5y9M2i4Yy8iu5dKvukSzia0Tvlg/+AuyZ6L0XpOM6Wfi7l1otYRBBvU4vUjuN
JIOPmFnw6wKRIDityFttKQuWox14rtVxUAQlevr0PamUT8jZHfrHXTjAQGWHaUx6ViNJWJ2cXNvj
gFPelVPdegNQyjR8fB/na10UHLHVtsq5L/BAQI3IA7UO7r6iXlmpbPsNOFhG6P20Wmnai80WJ6IF
MTe5ueq6ZMRAJN7J2K0oLNHGVGa8McugUm1N+WPHVjGu4jkt8LrkoloatAppu3D1xHKfKILUnRCo
kextYjmp9me/8pO/8fX+FhrhZByPem4uQsn9wGkJWcPVDZiGwbg4J9bBF/xgxABy6zY3nSRTLLEs
JXO6K1cH7Ya8s0mufmsLtcgA0NqAilEzIqY/fq/L/5npnYheIU8EjoI2lyS9PNIQS0+vOl0gvq5L
zpAPZScEBZVwxBScFdhSQlAeKGdnAK8h2l0O+oIFCN6lmuHKvn+jhR5ow+/1N9j6ueiRbrS3gR3A
a6ESkTLDggA6t/XAgPhZul09GmTHQ1KmjWpG+t66Kl1rq/lRu+lQkTsK8NJdio14Uii5IitHD1Iu
0Ump5IqWJ0CbtM0DdQPoUaCh4ByVsfhoQbmRlYx6VLBSST7Fs38ea3dFqf03ixCkP0kJlX5qHPaE
WSFUFmYpTzSgqopt842O7dKWpBqUsn2NnrFmkaGkmzVxce80iHk+GlVyYSp9GKhh+Hqg7Ukj7+3Z
ePTU5eyFn9CflPveQKmtAKySUylbuPPBdPz4OD/LMGKnUc/R6Ls4QvXda7YrO+ixnN7oc/E31yVm
Vo7P1RbkYgl8X/WPren5mPSmMFxJLxuGjD//IzUFo7yKcyUAqzq2N68hmkNj8svnofxMZrWrB+4Q
0wn7HMSr+iep0rQUtG+SdxJEvM5f1WJQ6X/rQdzVzqUmXyq9YyDziAvRNkle8u7fEFMmFn2CgoJW
90BO7saadeKmwVz+E1lRK7ZibkV16/StS+22DTAuTvb60Z4CYqIPlQHLVNqIwd7ye2cGchlUdhtL
rKUGQ/dAxdVIgmEMObHPZjPRoF32VezL9IFlgpQ2iSqz/x/mKtXt5q+++uOuNWZsPGvmTYYjd7ld
bpdIcCqO1OzQdTucYIIfv6RRUKu7W1BEPf+cxJzvjmHUdpmKJ7qyLGdgGWfH9z4d/uEwtMHuJzxv
UZyYbyB3iZyC95vHL1+NDEifwsBlNz1Z1w17qrunpYHltFbbyRJtSPTJ5gm4ivqIP8DyGEgPdgNL
K7/wiEcr4HWfXfXESbF+GHjp/HlAeXHl+ij6O+POiZ+mW47cheFsLGVV5Nqx4vTKl8WFkfQeKIVr
3wuM+U7YYGYiGbA3UJc+iSUkSis0Vf0zNI5ZjALbtNFwO/fT6CocVDfhoXghfNOq7RgJv2/jxkur
KWxZ4BC0PglhlcEuqtHxRSLDQHrKRHL891AhiCtc1itvmdxbji0OraBKinc9TMMt099bZUu3wlJf
1Mw8uOIu94Ks+pf9VZ7WT9mUar5oYUWrrS4WbktRIER+oh6zg6JKvMZdQEnA1+W42vmdhPWRhNdJ
tSXtS2/7bK7PcBDmPVnj5uw33EtP3eBV+GDoXuegYZiqCuqddrJd7UT1VOcCPDxjcGCHgIrK88b4
zQofn0iXk5mDak7Kx2MSMzB03fcky9lBv2UAGgQlhQC6MUEeJiVIjuABrLea/073kUgjqHBvLtJj
SO3tuln9shvQWTktBQSsBHvwLY7dBeUpUinniPMeeLvZ4roWQbBC/4HRD+S4Nsyj92R5klB7PnRg
WOOqV6PgIYgXQYMpq17JDdUZ1I9qIVACXgOjzjcQfgzM6vKYiZZQFAXMNUAyiCogWywP411xP4p7
2SCybhObuwZVkmk1A+wYEXaXE/nQTy1UiP5uIaQtJEZlAXcjq9gBIotpttfm/7A1WGsbmZePA7dP
rIk90WpD3V5Cs2bel+gMzIEwHRkROMKvr2bwIr2eaG7jw5DogbnIxMNAE/lT2d31Vhq1fvbL2iqw
iyk4ImojfACidgkshWITdWHjAEDZcaG/TBMctcqbPsz5B1rcPW9vhy1JRLAcdQA9BSPCpQVqe4b9
WvTJgTg/CAtigr7Hxw9TuqDBtJFj+5VUY1q/a03AKRGVFD86CYc/fMLNPy9veKa1huRZ4OQHE0mE
XoMjbO26idFkBxc/tpgoRSOydeWGeY06R/Heho8lt8P77wvvfukhe35DvcoT4NPpBX2tXLDQoB3i
fCTW/LWHEiKPk7z3hokuC1Zya5/nY9T0jELZ+VnHLvlgB42VsAHj8Hl8AJzFcX3HwelBUMh1hrtr
CsCMdl05X5Xq36p0eUFM6vPSRMyL87SabiKqTH/er++Knnw0Bn+9/A1DqusXq2zA1/R6yap5FjbT
GAr3aoDZJVY2bSR8aA7yH8a7oRwdiPgfGbJaz8HaVtl49RGLABfOfUBOMSwqkOYE47Xq8J3OEGxb
BQ7zHzCxstmNkt/Fb0Ll+WS3Xycz+oOSzUlNM+Lhr7vh1Zm9yfiyiUxq4CXGQzaYwb/POa9CJOHp
JSOvxXqSPPPFn5lF7K1zMLPohOYYOHhzPxD2JHUTzPCVpBRAMWH5lVvpxXzqvA8Fc/JaVOTy3uxn
ZeqmaIG30xt2aiA3+rdb1yhIHYgNtyc2eDuYpaLqosbkQAgu3NUEe1NQSqKv/joV6SNh+uL4BXta
c9vkaBDiQKSbLezR0gUvGXixMd2tSpOos4ZzxRDHG7U1juGCgAOB6sX9lGxc3yq4D/+b7A6MuU9q
dmNVunCvxOnxUeB1jjn+scxcKsQLT/o+ENa6Oh2hY2pMAOlnw8UCDxCaJ7QdyTD4hpRAFfInSfJf
vJ8lBdWevJgyDvV2MKyilT1aUfuht5KPtpBubRgjkTOESFPNu1wcNwulkWCnAvtXs76I0KIylSiN
89tYigK0tEI4xQPDH9m7yNTvSBKQMnmqeq+EIJ1f2DV/KHSiKKPBpY1KyZeIx7j/VwUv/VNPXiTa
8phRrkkpg2s/5HS0vQVR0GSxbNj5s/6JUiT2CawnAFwLKTlzk+EFgY6OQezXL4mx3FTt3bP/0Koi
Ugh/S8v4d3WbTXLCNOZ9HqsalYnPjSRh2wlC/y2LHnMALOqHl5ciJVuuOhXvNq0XGJ0xGSEWL8ru
mjtenioE4xqxD5j5tKumuL63t+8BYT+PlZtfibvDnHUN4bgHOuWKmPvf5oqTa9vAe4wZr+5CanI4
bAAva3NpTVSi+4SrDNLKzMlz94AZv8aQ6+kfCKRUBiZcV+FHQ1ng7dYZdf0qpIGYFdrWLtsxP0Sz
xSrUSr6gRz/HCOy8GjsAQf3znHIagrMarBhzj/j0EbZ4e3fnFH459O9it7DSjWOHNfZK65I+mw5Q
8twDJwL7W4XfcKjlivY/oAryi6C7MvyVxWKgyATwyQQQwZuYZj6NGXImSi6iu9y54sh8nGAqUUXw
F+T/4H2zUBI9nCp8d5654u26uV25L1au9wIqX2zSiDK7Qulew2tiULGaLv3tJVBI/jBDF2XVnnob
BKSBVN5qHaW22i5rytDjdm3l+7ORyKU2ocCNwNKp/ue4AKVEDuTHxqaN8za0ce9/DtiiNEoWEPGe
5nEkPjW23I9Cs9G5A6bwVUpeONaijY2RFcz13IhRot7Epj8r2TQyM5hC5bP+/dPz+CfW8OzfLr97
k9T70XBCrI7/58sKYgMIgmTWVGjMOHKWP24C3whb4Fx3b/Y3tdy+IHHgSI3cijJ/ZG+JalQu3g5k
rQ5S3WyBDVa3nzB/0iV6pbGxaZD4Nyr1d5i786GuJuw7ffW7lzOm2V3lR8OzSoliUr4VyboMp9dc
r6mOBC2T4Cg+CgKKyzF/OoIkHDTBLinTmc5KLpJIxUUZ6NuCmUOrKjEElcDuvJ9pAk8P79yQO9Q3
HgKIN8VcwaKvJu7VeHzVMz90UTe7y4tiO0A449W4FVGpSPufU4KAq4f/F6oPPWRbT8D1WKauVP+9
1+715ZOZk6sESw7AVDUw0319YaMk/85SI/lqbhbncgs6pI+vefxzHJFd55THMqGtcoIvFhpEm2hH
k0zyLX7vstdCyGcHjRiCHbJ7SGutv1E+mRN4sGhWAS79HcZgdxK+L2hdSgAWTg90YHFcPtOSUeUB
FQY0scIlbkMwWlATzXCxRk4B//VNHTW/H3qZObT0LrSlV+srr8PbvTd7xt6LZPQ1YCWd3zkA2iNf
S+/ChO2X5Vrz21cMv+CJ+dQYRPybY+QW5yY/bPDodYUBjBE66eAj5uVJzUWQsmnJ4IziLDkkvKBT
GVEETEduAhKuXTg/7qJVUAuNX/fkaadj6HiZ8j0HnzHAgE7vCHQQH/qjyybzO8bJx/YVi2SAICj0
/rxBbLapnutlp3zIUYJaKuhSMLTlfZthN0RByY1FZWGV2N4bIsZh3Hy/Z8o0T2qg/x3UphJU6f/a
C3gmM00DTfco79QnLNfHQ0hgcmdq0kYZts9uI0mE8m/IUDoAmbxLF1c00NSOkZMBiCpgpt7ZjXj3
2uv1hmLNHH5JCk68ZHq4BrPec84OfEa+iG88lI81YrmeKVO2FkJt8DwXuVS2M0F33TG3u2uPdAKg
XQcNMZn9AkjkJo3qIq8yGCIj+i/c6efLv0g1DFw1cHLzBBF5EuBk9MLsh7z8Nr/M/m8OI4LdOyir
4imKx3e4SZxac5uszQZ5bnjYCKmqaV0cl6CCRkAwqW8jUwcTVfAAFbZg5mR8wpsJYY/3X4kAijxp
inwuNE1le4yW5CZMvMObvHdzBbYZnQ73s7WeETftIA/X7Kj8GkLR4mFlsmA8MNEXKBffIb8IlYGY
B9qPBVMJkaoEyLGzwDgjCj1a3kFVjmJ6XTO5B1xroSj2QRVkFoXqgSZPRT1TVx+g2dmefcRXLOBB
jhLO8hT2fzGDnud9AQT80u9ziJGEtCxId7RHDEdVSldGuAgQlhV+7mRnAu6XjM5/Woibzc7NCTti
rjtjUphMQ4QWTn0FA4wjjp3uFoGjQG2TC3wkHc3Wdlz+baHWOL0ywdKHQTTo67tDsG9WBd4L5Oo+
/BElfqoLt2W+MxOQYdZjhxBb2gQBbnlAxr03BwRG3YyZvOlCids27eB2tDe25fThKHAdtejqOtNT
zHn/LSrNVyfKuRNrUo01NmsrdF+CKuZ0KNGAyhw0YxcgjUPcaaZ1ZYurnGYaLOUI5rnOzU5Ifmev
ZYu0F20INNtPBlR1wusWtHNGszJUIX5LhQPWHB7D6FkVl1a7fPY4SW6+Aa12qBnjRSbMIz36nhGN
u2b07jc/0PNsdz5nJIFDzBw3lXHt7VTRLtqWrizaoVcvJJyOuroQF9mmF/Dqq9volhOtYLTl5nlx
mjbN8axFTC1MK27sozu185TfTYgwMcCUxtMVbAS0Cr/Xb6H4AhFf1FKCtJHI6QdZjxZIPNVPbwsM
MdKPdXGEJef+gCMuHMfsioqZc+fR/16hmeWCDAfBMnGZmiC4bwx/mFFT49rp7R3xcSULS06ihz8B
rVjKCpBa0zMpxbJjUwI8pFQQx7MMUWe8bKaKUm6vjPUxkHIO2L9FGV3kdtz2w5QXMavFYQ1z1BeH
z0318plwVRW3LkG7XcqSX3N0WbDs7Y9rO+B4sZiGwLnotBG6K8fuKDqnglNrva4GNmDi/pInFaMl
QQYoV91pucHQkle2UyM1gSIpeCxyZL8CQFZN1DyYxi+zceSBmL4avnm6TJhBB7TAJB6b8/srL1S1
Cc+eWBa7wcPbrtloryc4I+xcvKtZiHpxcXgpIWAaIUXnnwemB6+QP2ANkMz9Ti5F5j2rb/LtQVi3
eNP1kK77rsYLW0Vp9GqcgWzDxMr/xSa4ft/RScv1v8/bTNdmegicRNbnX6ZCh/dxjccOMcFPNAud
6BkVyHYHov2monn0elaBopoStJcvNlZ6XDRWSiEmIDg8fDARmVrXB56TCr+5kzyDRP19OYCpSUAl
/4DpbmSf/l8Y8WinXkGwzdNS0Nut57Wn5HM3eyqWGB11gDDNzQsk8dhEzLq2XGgaUIgdVKUuhuvb
baFvSm6vSyREl1KqLMYEUj9fU5PcpltAH7tcJi0f3rf9+SkakM9ZJp6ZKe2zIsaw4xq9+yarSPX+
tHN69OUw7ZrFmsihjjAhtWiimCYEGzo4xjtP3lCuFYHK/OzPfcKZtBDEGVGER7QqFSD66Ag+PA5C
8q5jJojXBQDi2MoxOLjQ9XRSXrJAUx6T0IVQossET2gWSKD6g10x1ZpeXhiG+gELprfhKBGiSfoz
DE5kuhMUv5gWL3NpTmR+hD2WB2QwTGu6Kdw70TcmWz7KIdsR27Gjl1moNZwIhpnimcXX1zR3NTAW
hck4o7aAh0bxyYLYTgkdjIKTxnkPoBpUNml9ARDZW46meCI5f+T8OQMQcGlIoPCQoJqx4uNoRs+Y
EJQSSm4shtnhtYlZALmaDvDgr4HshHoF0tU893iveoEocGO0II5gUI2OGD303WgYGjntulwJVLNd
/BgcreiR5VRg6t3dIylkFcnOce4jAPEVWdrGrb0+gOgBlwK9L135sSba+c1VBeoXf8xaf6N16wr0
h8+wLnu0bNAUFTY5jDxBwHL9Q2d+Z+Vc7BoyKL6ITIE1bqeuLBQCKKi/ALVefXlBD4OmtT1QrTSg
4xljOlOUFJpxHdtA/guGOBOz4rRvsDkHczY1kHprn+o711KQLZyjEx02Is872YbkmiF1+gfBIf9t
CspYm0guKOYFT1zLkjGilXFytpN/8GqRh1FODCfomibl1e5NCrS86whVS30gxQlLzNKMTCewPTQC
zilS3WBhXMPbiouswK4+Crff43OKzaWTyisgPdOtCVHqlXEGjkIbHb/0ZOCZCYcJ+5hQHGr5kR3S
1T63HKqJxWuJek3c4FfG/5x4i+eJFgo5aBiWbHbHs8dpcHAtE9n6eeKGehZ2vntP2Cv+HvAKoQ/j
PuH2oabqF1DZFnyaIA4k36qfJ/kh5+y59thEYZFGER0vs9A5LdzfaQv65VW37Spq2islHKHrQBk7
kXDiWEW/0I9dyP39QVwLOLbXALSjtzISTWIZwg2TD3Yn0F/0licUfdQrfgrawp7AN3BCMnZt/fjK
7Lx7VYFclLjFcYV6h1FL4TLecDiE4kCeKuTuQaGyxn5ZCaDlMRRKBAKJI8BUjf3X5TuQsDTNiBbU
RJmO4qScWgOGqhiAI3cBEJdZPI5XzdyYDyNpbevE9zbVy69Plm+b0RZqioMrN7oAj7rInqqxgiKN
yBBqpXEIW5n6QdNXzAcM7Tb9UEgoHZh5QyObBhuCtOplMf1l6S1TIFvE1xdcvAFFCgLColWFSKrg
uV6rhZmsZo7eqczNqSGBxie8uAJ8W6kW+YI3mRvZe+SCTpPULvyW8OQJL1StIZCXXKWp4YGyYnOm
6k60gBmjd60qkyO+Typ74apZEyM/8LI6wT7Jl8Hr/ggYA4DLt4GT3qJy/UvZVhXrz25ikNiAolmY
AzVJsJdFTD0YtVtMt4rfcNrJxVRZSh0om+DJ13e66JITY77/27vBzif825FBbLSqzcV5J9noXDeu
M/15UE2ivw/rlH7Bm6KJgq62RqF4XIfUf5WpztGPdESwSOuhoW/9+aWAUIt1hWo7PxRyhg8NSdlE
r2UHvSn+p3dbttk10WWftv0OnD94f6rRYM0sE6YsfP60P5UTHqek/QbZJJJeIPzmhmP7iseHWqAF
RnoAoPxe34n0G5vs+5WO67mynd7kGTmXohh+AW+srDDW5WI/2okGPUEzRIlqKrs4AigecWrx0Dkm
lnVSdRNwbdjqyUSHrLzwKXn2WJnss8M/dPJbWxgjQKwHqZrbaXSXsmQIW7wafz7nQEwcx2OGv07u
47xDJ4mJVDC2N6EiLbeW7YWoJn1P4ycT7x86BOxLW7lyuZzfxLUaGfJrgsy5hCm2MFBgBAhKC/AZ
+O1/0jj1RHjW+5nBCgBLRPHrlwpbsnOocNeZ2nBncsmm++tsxDGlZqGzt7ImbppoiHefi5YvZuNn
CAi8XKEuRiFdEyLfU7lhgyye2wHGGepPB8gunBTs3TGfENAx4Ibcq9lFv7WYcBrgE5tcYlt57iS8
eNMOXwA3hqLmaHo2c9XHU/OoyDVuRuXoa95msXJu+qXX2p2g/K/c4ljAsVhN6L2INh992nA4nJzx
G9BK/+cz6F/7uLjkrt91Ec1z3GXgbyY0Ah4Z7Abe9ILMJxQkOPk96NP4DmrVp9SmzVvweni9ui+9
yeO5kiqy6hsVlIKkfDoDzzoYhvDaNm+gP5xIy1bFTxbB/P7nWmGzvzrOCL/Gb2XGNPRrYG6cKAaS
VoiZKeDlWejtQoGebtsW1ITpr1Ogy8czPqVD1gVZJPnGoAFA08Z05JXNL/oge3Tdttb2fQOQBS2G
YMMTBrR5FmQHbKY4Ew7gZIXFeJPzZO5oDqmrnK5XKKq2FqpRlE2T3VVjPw7+J7ZpmLiJiKMnm5Eq
ehIRamnhnb49uC8NLd+h7ADcya0mBd4u9LIA6wQNXaY26XAP/XzHBxw6saGoxKBYFED//zh2tsiJ
HfWuQceKvJ3NLTvi8BMn5rQaeVL8Tajn3MCLhfovBI72dACvELk81hGPwJ0FTAAjhTytYl0WQHDV
bOIz2pyRoCM+iCcqar/g/DBJn+5TTipbQuO6iAPELKoqrZVwUIukCbODrO4dtfdrkk5uAsEEOnCB
Ll4QeXGiQQ3KsLzRnZUJK/2OrbkVQ2RW3nwP4yNIXHfw39I8Rnhz1kQixF0K4bVdmj+JiA1QcdUD
ywtVzHCY1SjFRhQGlEr6yGAU0IZzuckzqQpfdaFD/Ea2L7KE4dPpsS7xeYxV7BrpWA5CRpbSPKP3
FF5vGIoseaIAj6Y+JNdprn9tUKu7WNRYQvG2Jiqi/CmhMNBiAVJRubf0lY2+uyZ+7eSBOg8xECUS
KjkqGXh3pvwsNw2+GzAGHVSvnbJfLTmt0KO1NiNZ22JtxtOSXAE4698UhELP+GWq1zxBeyZprMSt
cr9Dx2rLJxl0mQZWnONonZGu5R+V6zEQQ+7Qy7YKEV3FTsY4MsinXBDuBdZQQG7xYzxwpbedbTFK
ZyAdoh30qJ93DZYt9TSaxinP8iRWpSlGQqPOIGPNZ1AxUnOcq8myJGS4RxE3xY7Q6oP9HdHa02wF
G6X5nU7+hV03nzd9fVZZXH8xEYaTLsV8dY8R5zfFj8B5990xzyfzwaAgp9V/YyW4xRBXroAL+bgf
k30fstjwg1EHUduG6QU6gqxzH24WwUwZ66GHhVQP/yY6EFSJo2vizjwyxJZD1Qu0r0XZYDQKFs2k
uWg5psvw5Hge9XikUrfEVxr4HKlJN8Txvzw+7ovk1rEblqkgmH3ty8UFHb9/MySnzy9K+BgmRajP
UDn6i7/pWSvLClP0SM7O/Mh6wolQevia4xs87zgiqWSkgRi35MVtKh9VxngNIDTtvGB+O5di6vUD
WpIDqSLhDRoQn2CZD0LeINXhU6pIIRJibxtBo8c1ooRj04zOmj/z+UoOWLUK6pTuF+oSIlIfWCYz
5amif1MjzQmCAXjZJK9zvkWIuJXuAouocrSH8gtYhiHweToYVaCaXoswpYyTsehUCSEtapXQjd58
A8/EpJ/Vq5SbabzwxPLPrrPCg767TszdjpF89Dyc8eX9wkQkfhGuXWRewE+4efCx0MabYxI9IXW+
4UxkFjxVzz1eqMn6JrAOqv0U6bPOjmVb6CFBqE4gp02lQGCL8W444VmBhlWGwXn223tbooZTNRi3
qBuJNst4Go8DjjRF7A0agYBMiws79rtWw+HyFvCxw3c65cxdLxHXrvLT+hVqCps8LP8kRisz9L0G
ObokxpIQ6WsFQqztmtx9AXKelzVu7QP4YSAqo6D89GLxLNSuoLwImI/AIsBJ278GmztOQgxtsdDo
wQc310Vx7wD7g0+egZSv+P+8KaxkCiy92CV4rIeAgXRr1CgS1JoL1Dpz4onszV7RI2uSgCALGzSR
0NWvWBnA/nUlZV3jlUUziLRhcKaTL29xfGOPsFec6ea0KebMJX7ChB1iYnqVgHVZHIDM36jb4CDb
aUheQNi6FV2QevVGuLbOHEzfjJcX33C6vbnkeXx2lqg/nHr/WfGIhVfbkdAycQqQbLi7McQcFPzM
f0e4WonqTIz3QnaafzwO2SMeXBZI5Zi5wCTUlQ4OcXcBl+khwICQ/FJleQXnXXyPmoJIK2XXAPXO
zMfV3xVtxdtZYyAgltWoxsIaQIU6+mjWikJvo/kYaV1SfQ1SUVx35o1Te2RhV7NPZv7ri2Guuqaa
cXSqVh2BQs4vIZbM4y6LN+Hrghkb+TfwaibWBLMsCuvT6rQnIBQ8O03GQQN68SHtTk4WxId+W1ej
1g/oiD53xfxNEgYDLIXWm9poVjXL3f+uLA5iA/dwD/1nNKodBd02U5HmJ4wOo5a1/hhmzAztoxoV
rnxoctzF8gGhhj4vJbzWEhdxjLvSNPMSmL3F7IXOvKVpDLvk2pW5+/mMtLhpPuFzA+TJG0i30PVT
DGEsx/xV7CCC9U+BLfmrgD/wJ7z4d+5jCJlAtJLm9lEj4NzD04zxX5mD5yhxMLBjkze3dpubNWDs
PPJMLYesgmm5QxfHH6agMwWudF+h44xlAHA4Z4CLaL/RsO2wOQIJy0pTw7NDqhxNoA1TakgJ0TgY
tejXLw4Bb1+cliA/GLyf5NKaeaW+vg4r6lsv4Dvujf756CtmcrMoFpFHWgBeNwiL2SvebNF1IssL
8avztjWKDfmHscOjXLDurPWcdnaL56iD3AVVXl3FLeVBITHPqmcgXBaLrla25vE7Wimh4TtMnMqV
aOJXbhsLGmF4DpyfJe743IEgv/mKk1YbgjuKLisnbIs5T2oXZZgV5Rti658PYixal0TQfjX30Qrb
FpjLlvsDKjBrxkRN+xIfXchkTcfNjoU5eNAJgGrgzWajnN2Ss58k5UFCGKIiCQngNMb1sOilCOzv
M/WBWUKkT68tXxZzgDBiFgh/pgoF/m/+5WdhV+mgPv2AjEAOSqrFeV8WO5tgTcYwqsFOzgETilZQ
ja7qJ2Zi6JW2H4Fds71lgz9nhJVk72QB87nJrvoW4h66PD84tIjMZH6rzZeA8M29iL+xpIgpSd3t
vTSjHoamjOLZsFUy2J0g7o8YsVQ8x3WnbT7jh4rwKy2+Hl7giGKKCeO1hE4Cg/rGBzoreyOtEvYF
VeGT8bGDEXR3Hh/n7Qtv91pgtlr43s5fcwDcvzFnqXFj3R1KXhIoc/lHNDqEfbX5fDUQqhH+I31/
w3Batk6u125j86Yf3Rtzh57yA3XewaiFAnmETVfFMk3y93iNk2f5cX0radJZA2CWIUF7S9asWdSC
sSH8eP/+0yRGQ5MLdplM7j8b7bWUqgaz58EJKVS9MPlzLFu4JhOq0wBHlz6bqduv35F25sV+RTnT
+befA3f2Gy2tasHoSZJMK7UzPyLQOuRYeu+PyihwDUyWpEome1ici+fKOpwBToFikXAJU4R+g7uZ
aMm29i8E30UeMOTmJQFlXgcv1fTt4CmkAsMy/1C6G0XFEvobOHMaPPJxXEnsgRcZbL7DkQEIRiJF
L09jzeUuSiFyGB2QeezFDyoGsoOwSf06phlOOJKwdQ9OYMvwKskcwlH3XPrmY7W+aqyjXtO0phWK
+LoSIzrctDurya5y8S3VNSnv/rZd6GjRVIQMzCgCt0Q/3RwHMqUphYmFt3lZXVKqb1Yy0PJdFqxe
Omqn/bnRJwH7PeympmPPBZLrq89TXQDw1PFoW29E5lg2NucR+o2tgDlIibKv0kUfBzFwlVwC/AIU
isaBa2sDTO8q0m+C8H22khe5fUATQoUY8sZAQa1Bf/Tfpy246s05aj89K2QKH1phhdyWtrI2IdL8
viYBSRaFZjrYHQC6wKyUe1VsdCWkyJFSZgk6wedOLeSxD654tmtdPJQOZL05QqzQ30T0fYqrLlra
/CO5XymH8o85xATNSkMQZ3tPgoIyMDqAFoIx15keCKGWpSglV1fqeIAJYObgNxLBE7xHO0Y/4VaS
dg+UgXjkRTlOhpPrUHG7o6e9I/KWP8QeVb/xFXaK9N9sTOHJhDRz0T1bLmZdiSmiRlwXYQ6onGv/
3DP1JOKMRuZcJUnd5ssxIR+QBYp39C2eBeBBNVTfLG9B3hI+tN/dYaWO/hKOD83TnQAgCE/D3iIQ
dmZvHBGaLEn5LaEhBnURoLieZCCvjXDDVlSCopp2zkZpxBriTopBTOSXg1ig3/ahhplJ+epn6HbT
KNPk8Py3FUV1YIlTeUM5P20id566/pdNMBGpLaE8FFK4H8i23/kAJwws/LyYy/D7/XcVdsNDobsf
N/XAWpk7SLHfAbSj93dNpI9tBUo/WduAlpSpCQHDKTmlNOjeG+zOwKrhLsoS9iYSqDFRA8escvS+
oRjPYQSUKrWOGI9j0zGlzdqtPLwk289eJq/STb85ZquSEHD2ndH0Tb33uAgQ2aoz8WJ/QhflVjto
2F3lnXYit+PcePVSA/sChfj7yEin+yCs3/89+kesHCDmp69Z4XusfdbOO+WeBXKQdrmuu+9Yng5Z
1HJjoo5E4xT+zWedGasP7Bo03cjrCmgZFP84r/A1vYMnPnzHClGQWjcl/q6fFS721oP+0y2yJqhS
+udbNlrfthBXSZD+JT6jDG0fKn8Bk8sV4xi4W9YdK/6RBDHldkzc9gBaae0nl/XhpbZVl7KS2F9g
c7Lg/10DzB+UAhT5E+WfrZJhR2s7dk46+N/kRjH5IPr1u30Ikqf+Qs6age1J9q+wUBP/Tmd/hNvA
qrvfJh47OWA1Kxxr6W2xLGP0KYbk+gIMVjmFixNiALx1Yb0JnbzJIowEAVbTU8yRAZovzfwJyMiQ
maXDzW8+OtdBctc89CyyCIsQ+DmV3JmtlEyegxMZKQodM3nqmjmd/pkr4iUY0pxS548RNUkvkQUl
wAjxzRGjGn8wC4yMSDoTPRKpiMIg6t7YhFgKvwP4nphWTGk24V6RVtMPu8yduObFDgN9Oh+lTncI
rBu35+cuLIHo1TpvryWyEZAVm0v9pzXIKUmQISldR4wIbqBCjpACL0ij5stuZrS0WUesRSbQp2qG
fmow+UeSYNSV+In0fnAhPYmfo/H8qoGikXT+qEYxzRQ2WbgRVY+vSH/NZsaW115Ndm2dwO/Vhnzh
K5uVVzrycSyru7U4XQoBC4zu2XjLeHmCCshIPHiWorOGe1na/Va9LZjLoWAYbbcR8QZgCFyHxgNN
9N+eJz0gSY2B7GYVvkGsoiVrdIV87vpmeuAlUXPgtx9VBjaMkVdbsPsIp2KhZ6Jc/6+XdvjKNoEr
Yh5RuEuT1k0qpqPmYzX+S+k5313Ut02HONMG9akck8F+svoXwoFqzO0PPQph29Zp2gUxc7wP0zeD
0lMkDeOhsGzLGp5oOBVOXsFQm3ELcoYdqUe6HX9z+6T394hp1BD82LOL4O4cMFEfdWhZvu0kruWo
lX0SCvwbLjCcBKsuK/WPnTmE57PzbvWGMkX78PDk2vbALxmGK+fINACv/fmtenduN0Mqo4PAgmOb
1nbVWQyQyE3MnsIR3y7QusvYuGzXl8ypRqx6rs32ys2GVr8noBcA9fitXC0TxTtvNzRqqzuXDW76
2BJ5DGnRDAPl4+WCmkhhWWJHUF4sGhwdNKLF1//NaSRe/qsSmg2LeRljMBQ2D00bMOjQHCM0U2JI
MSQzHhGTD8VHZSbCgyy2fdGTdNyDAScT4rwN580lAv5V9mJZhllgLHc8XfCP6FPSQiyWcYJPD03/
8VUEy9d4amK3Ca+r//w5HZaN4WNyduY1cjkybJ5A9zvv3nuH0EMd76kIub1WP+FxQEM9KwFhOEml
5mhF7u/dlnvRsQOl7Y0cjWEoBiTP2xo8pPanhlt83B+pdTUlpJZAQr1wZ3tg6jA8Ik//U/Ppp46+
XZZex7Cu5+Dq3YhBSEMdXuNjVYjDBimgIgTFwLSPb2TULAng/p+sciF5URyPUOMsBTuIs+ILI+F6
bxANSVjz0Bh/1TmsHjKtZyqtZEku+m0DTLd+i9wFaHGPkS/YITx9aAmI5kY9kBbj11I1pPbnXZfO
gRyod91KUuj3MaW4e3wj9NKU2BWTeBktndent3f04PpRzJvmefZd2uhcvPljCV6I0/0kodaloTXW
G0i6sbKLv9MhT12ycwaZN/MO2I4MblBHvQPRpFeNnNRgxUN6xR/KLbehsB4lSxNTQNrBp1NqQs31
KDlUfewTWi4GvHRbVwpmMPsM9Gi8Ju8+auGrGrEaiROrwp+JKJiFemg3jWMFE2K3Scc49Ahh2Uhh
kovej+iTWDJS4vB7O4RQ3dYbyt3WvkTJ8e0ghzkJw3iyyKhxjx8B1ZcohOQRdqxfjB05cWFxGclU
C+VRj3xBt6loe9BtbdpQOKekV343bIMu3/rQhANmu6dPKboV0giZ7iC2I5gzIMGuSmkXOsFqZHyp
OdlIlydqtzaouWmUCfDK5b8ud0X3kYKtbAY8bGS9e0mzZq1Xjg56hu4sbKbAhoNZTL3KysERZX+1
th4jV61A8a3hcEtpVBMh0xCxWkaBdXsFzUzIoKZ+2fj+CfAFn13bn0nl2RR6Hzg/dTzm3s2bN6Ml
JKSg/pvKHT1kiD51EV4+/yTLk8PFItJCT6DT0D+3cZgtcs2/JdN76WQExYuhrHISzIOQAaDWTq0M
qOAniY/A1FiEqVAYkx7aaPvWIHQ2rF0PbyEt5MDMSOPg04Cy8GvxUo/FRkinTbK58iYEfxIiaTg7
XHl95GtTbDq9PgQ4mx+Ef9cm/N66C+UeaZFbVwDFalB4ADNmNKvaPHiVh+BumEf0MgP8+14MUAHs
C+CAfNYP23VRnhnnmgG/GSd6ICkeXoQQ+rwMfLSazFkC4iEV7NyulKShD53W51c2ffKsv/WfiGtC
Lj6HdENJIBFGXUbTs3CQSJQcaTNKVIdKvF9tBQmKTAdZgX9JbXEu/YCoZS42PDPcbCREBjJ0pwP7
SNdGQbqRx9i/ud2r0nLtytpuNTyXz6anRJnYiDh5nJ1BIqB0IJDijwxecozrQD6XWak9WUg9CKo+
UiXXEhcJRUI9/0TDxAhFhD35KgN+ExoPCQAgIMH+F/xKvwuGGJ8kgQXbdfhOyK4f3ryH/OMN1dIY
Mw9/Y+S1+FDVXr98IprpJJJWk6XSbLxWyEjs0EJzSG2nrKeTeK+SvmZKQQyDyQAZqFLfLd73DsDt
3oRU1m2zkRyNsj/7jUR67Y9PYzw2vwCHm3qoSrPr9cMTXLn6/hCWlDRF9oHK1vACMEh83a1sBMBI
RsJ0mFQqPI4VdU0CFUFAL6bzWWq0yBhPzDSYoBvaLV2ZGKE+/LWFj+2b3S4807Fs1MKqNQtZPCSt
+roliIrWMPDD33mQnO5whno6zVVzuNE135LV3xLGYpPP+OlOVC+3lZb2gSwL9aLo1ZJ8wfwRR+W3
cgiP3L6/hbRPezTgl1S8869IXjjodg9WDFbJz5F8sYL6dCHAaxwyYUq3Ty066j7qtCBAte9aiwnr
Ez+wCIhMP/ag0lA53gx8DDwUp5XchlD1DqwruJCTK8pL7CT93ynCkgJT5w6LeOXhHsSxxGT9EHjo
8XQw3ZZGot6egvre2+R+rX1ANIHIT/Ul5osE1jXZ1JIrHhzMCO+0uiXjP16Jej4TjIN7/MUjnu9D
qJamDp3XqKeoJ65+lkMAeL+RhyyhEnzvyTiCCf3c/1d21c21HYvgALfFXisUmA3SJLIIVDin/13f
ch7gPbflwVc7j/Hi/cZ0tFmr5r0Q7//xZ0mCvnH2HqAf/HXm4M/Xcek69K3GTIlruZyjtB3PY9Lx
TlnOEo/o8Z97DLuuDlwNLjucFLmnHaMcIU9vtehILT46QvdVLOc0oCuHauiCf/n1cyW+1XPM8i8G
IRtEFXg6AIKTW67jb8BIUKtTS5OyX8ieUkbPYm8cBZDHrwQaFdPHacL10TVl13m7zDeZehRuEsbd
CHgpdoi4lrDpv4Iw606buKbvMyvXKdSxpX6KO8ZU0wGF3N9uDsUC1ApEeUiy89Qn2oYJsBP2UkAD
h2k/1I68EqNZX3MlW7vOUGzo5PUj/MCQuPWNKhkIXD4FDXQA2vhHCClQ/EYp16y//J4onSni92aV
hMEcN/7eY/SBQEROz+pYyOmZB4wmF9014mYgNzC53N8l7PpdrVZ3wK45gPc0+CzuQWxSrq9663td
xFFHk6EH0vqdl/FAyv6g7rvrncfP+OVddDKx/Tw/hRQkcydx5KzaMoJrgEeR/hE8DEOnU5Cjxs4N
Y1K88XSc5Zk68GNR6eOAfQGwNvaxBko/XEQtHZx2dMyuYVlSGS9abydE+OcBDrli3mik+sIVBFZ7
mK5ZxMJtBJQ0YhS5LpDiKedE+J55XJNOR6S2M1mdPT0/QXpmOhiT0+KU7vNWqhB8nQm2PFZ4IgIw
Yyl7plaVG+oyZFCX9+Fi4Ie+2omOOdiRv0hI2T0ZbdJhwyODRYiomBDxwMQNOAWxI86qlUAxFLaU
L2bwnfr4TWAA7GLghs27T6I7AvI5xR8yoTEQ3WM/2rOl+ra9CngfatNaUd5kZnmL9FQtCb9dC+bh
NGEAe/uRIi+Dn83HXpktTsGnzHUfgOTiZcnPHkfOyZugLwK4C/uuMCMHsEPIQrixcRUd7lvi5rTj
N0qPnA/298vxHAmbuhtRH/Tl2HP1pM+N9ilOFGNe4o4ZhSl+THOc/V6wIa92LJrr7Sa1GiRYAjLm
vwuFun6roOKtVvfv88OONFL4XilJPEnvEYfjeoPrBAORhJ7owt4tOPWqlmCT8UDYxeB4XJcX3eY/
6o/eTAljdM7HCCRqD0Wox2Hrq4H8M/wMsWWd6y7m9uVKF7xQp4UG3o9TUr6QsS+cY1GWLIIXc4xK
E7MxceKDtgI654nCbQQQmbotaMLuoB8PEebmGBnkFlxAaX4DSyOVZnAeHyAJggkZIDMoA/kuSZzj
yKjxB9W7iuEF6Y0rz1juv1Hel5/3XhjpDEqjVZGeim99Jsf4wnjfxEcSvheOpzTeuL9DIJO+TY/Z
S9h1JbkGBK69rjgahZcgp3BRvcIcczcdzQUXPe/HRN63nRbgTos/qpkx/P/KDAwj4LhnF42/JmSs
A5G6QkS6/+k6gWChmiIwBrbLSam+Pr0xClLWS1X4GBn/8YUb8NpnN9PzRyOqIOJlGued0DU6efPK
8ZMtB5t1pWnRySh1GScYfTAHfl1XTbSArfMuES3LgGupKQLnI+RnVNlTbSILK58vTEZMEVDjSd72
divvgt2xdZeCGn3ojljxw7pncYWKVW2CFGyrrZLnDeWGg6JveJHEX+dNErKbN/HqIhdTWsb1bYFp
b/ccxCCqm5Rv1Q/s+KgHRmkz/HV0CzJm1liGuUSi5oLOBn3uhq1Hd5F9CNqmb9+CnY0Q9/aFPkdK
YCcHp0r5KCjM9AlOfTfv4VJGMleBaGt2uJ7ogp3UcHZe0wArxC6w0E1a9H2jLTvZCDBc/ltWOAru
UY/+dJN5scjeuOZnkBkfa2lO+/PaMDGhfkadeJdLvZ6L4JPcGDbho3mHBasil1s9T+krlTRl50wf
TmAhQjK4/c7HyBwd68EG1FAjvwM/llrIw8VcbL7i+UBRfYMOMV00+EP+SgmtVUKpZTf1me3irPPP
BmPlBZPYxyp4TPGvIfMtbuEtX2Ul7WfpjOKHUmS/NPV7gUzzsYSAjAW2a6aBTS0QwZRDxJhdopSj
lQVvBaJSfMyDOXGdg3vaaGcVltbLUA/Eqk/UtA8A/qG5+WmB2OpRc4p5wVra1ZBnjdej05AZbdAO
7Q8CFAy50qg/kP3BQtPXgkd7qQ3o10r6qXh0pQI5FuMdAJGKxftM7G1RcMdyee3Wv/mdwreeJEB9
W9ZJVYuvmw/DjMRgPPlKDVV3CnhJo98g2fipEst9ZT5JdnolEMfeGW1WlXlJGDNShfGQquhQcYWa
Poedjwx+dux+ds3eP2dk4ojKAUPxC3mYbXqyg3sSuftWFfskaiDbEsgaty/Swbt+jiWmc2v8ZW3f
yU+kYHj0w8lHec8PbhBrlyAxMjWFjYyfqcmORMR4Gc45P1OOh33CUrDrUrdEPP9ECeh72aFKIjD/
KuQUnjYwzF6USVXXx2oninmZX0UQhkcEbkT/jukUpp2RCjVvNpkpqktRJpZF703L89p/p1g0ny85
Ykya/ElbG3FU24cJWWjpBJeS53IZtR2cSJZDn2DZv+YrZ+kRniX3cWN4uYKOvFb4LWZo14FbClmC
td1CQxFRZLKVcar8dDE1FzouRzs4dh3NpMkmJmaAzWdZ4jaYwFA4yiPf8r7tx+BgAbSYeJgOuv4B
Py4qfwlMWqAfGp3FVcfOnxQxGL2VNjporpZYENJzqMHn/HUOJHBG9VSGfAWYFoVa1U7OMyrNLA2D
0G87TLLy3d/eh5HA1Rp2QMLDN3+BqR0t4A2+if12AVYzNay1pFAcor250SP44YGU68dVO+/rESyU
ByTwtT/zxb99c1TYENtwbCWGrqhEz8ALCIxI97Di+Rn5uM/har55d5GPWmScWAchEMlVMB4OxwVC
CzbHb9Hi6xyfLE8nUpnnQ4B8oq6kYoSAeN8zMAM2Uw5bGzB178sNuzV3tt3zJn0Z/L3YVmJWBYt9
d7TbkQQbw67N39CvFC8javjydXjxp9M5vWoHyHJwh1CSmc2CR01qSK/KdhDXq3WX8xrkPfyExGrC
RCH2m/74ZP2h/k+PzV3BPQqStC3z4ms7I0/cXCxevFx3q3Gt4CrudaNihQ3JtNniVJi8Jjl3iwt+
E3epi7mmZh9cL7VEtanSUPUSkfbDQPpWwmariW/Snb/oznqEQqQgi1toYKn4IL9sXah1DkH0WzlK
PKSY8j5y9KcdzMibFsCqTyGBnI+5Xsmx8Yfkvwq+RZBNYS46jzr8Mlwq/hmZLPg43A34zaxoqXLn
MsnKDJAng//2l/q7l+ChjQarRzbn4xZRlRW1F2hVd3JqFUMo+miFeY/PrpujYXL1OlRhSomESu95
uxiGjrpRig8W+tGzFBSA+/GP5TUhAsrUjMtXI6ROLntYM4Z6z05aM+jPvsE0bwLnQw96Md40bcG6
6B/XxefXs2C8R/e51fOQyVOSs0eW8aULoWZn1TCS3gQQZEdadP7v0rrO9mWuw6CxsbzcvKKmEL4c
Z+N3kaKnde5u7cdLsT9oP/8N4KMCnHUl2dVodHPac2eIBiyUXlUFPWIF6SHbgmsvghQaVQRIM4uo
w4X30Q/IsZk9lhOco29K9E9T3SHVNY8cyK0pcYufEa1V+fPlYUR7X/Y2FaXk3W4B/PyKGLwaGo2o
RcQW2Kn21X/9ri5MDMKIr6tQ+ZCLTCMomotIFjJuXlUqXXb4GXQVKEOSSZNgP8+p77rUWal/0b7t
HKXZWA38ubLhTfBJz0CQCU0qq7fr+KoZrgmUQ+nlUgSCA+OJuOIbZb+8+Bjn+ObzPz7gWJ3oI4Y0
D4FHlHYeZwcgElAEwbXpD7m2KJFMIefbTdn99Fgjp/7vdVbzfkS5bZrI5ANlktRdfnYHxBZw1KrA
Y5j5uVLPYfAayCuFVwbXb7R2vDvw5kC0i6kNcttFW1nWQzUYZjv3rTDwQ5KR1IY3+7sHAjs2Uy7/
HQGh1pK0mfppQLc8J87ZqlUmXzt14vkv47YFjzFAWEtGZ3HIlwfxx/7P4kt1mNhdCyMkNlnV+cRS
vlTrEwDnZkKSXOCyNEy7gsHWa2yJEKcPhIHNGJwyxJfvvwLYErKNcVtm08ixQgqQKcEp2MoH4z3G
gGXKi7cep++hhlmgOrvHLPdqnLDYVdCsQzc7c1CSgSCI0mdDBaESzycuYgJ7ZZxi3QgutKz970q/
AuTNDEQ7pVL5W2cp9oJy+4YwrFsP+17cEGBN/3dyGfg0CGV9z/cxYLQ+hHJdwwn2Uhv5y5ke/g7u
gOULbnGJE9M9M+Q9rqpAKT4eZVFdHIaYPBMyjf49s30ofSfjlB//f+CS0PGvJKHJSsUtaeuvluSh
laDkm8n7QpRFsZYnimTpgDB6y8GUGluuJSpl4BlWOES6Tlmwy0dEx2XcxFpy0jGwbhl7K5qybNTY
lmnVzHX438dDtcRERLr+IUyIyLDWRqoeyS7b1MjmnBvITxe4OkkxMUl1VFofP7UAWmAxEqUU4dfc
DoGph8neJstf2HkbFASpjxRVche5wfvmeI9RLKcl002+yvXXEJrsDWAA3CcIAmQ0jiBQBTX4o1TH
kDqQ+Kw/YcUyLrJWnKq4l/0PkVAVzVaaeUV5TQdGHFMbq1QPPk6jgU1p3+63u/yLha0OD+wAAV/k
FzwQ1Of5j9GipI1/miiHZRhUutCN6BO548LR6cs4O+ajYXHkqktGR3rRuRhea5HzzgkNuanxYxDy
gJVOTA9QI4wwO4LfiuPP06USGgwLywZS7wsjBuI8UWBfSBOY/8685ff8G8w0GvFHdvGVeGvE9eBr
Frrj/pQG7lMd4bdgobe3ZByKxfA+N3A1F0mIxezDUhe6Xfd4fJ4yMvyb+OcAFwJg0j2Kn+IF59Up
Tc9piIBGTVvKiA/MiHfUrR7sRTDzxETJRDC/aOl/GE9N5EIpdA3UztFTA3zIBFD/960mH/BdEQ9w
ZdO+KgJtR/Y6VgiY9vhHbLkmi1Ak1Eg3cetijQSTkqlxBLhlNBztwg+B4Gcp8IkSEoSnbb9poqvB
9qehy4zCp9tJdhWSXiNgyRy9ykGyNyjbzYNWRPCv4OB4wZ80pW0nCYmRJycp3i5nSFB7HGCBNoYU
/FVsD/OBtKixWuct1t6JrQPUm+Vu9L+YBbMRddN6wANStI4zEbNLwEQsX8FV5sVP9jHuY8mKa4vf
QDu/2Qd5BOO/DPVWnbFoBcnkVGwyXrHsDQRh23xgZ/0J7Wc6MsbDJ8cGfvtcdSF5fELdAaSQB7Ns
lnRnGOjDDI/Dt3Us9PBnbcdI8NwBa3u9krOmZDXi2Ynn/iVPV3hhAwtNzstFIaOlrKzEizokmdNi
aKWG20vEO0dDIbYf5D5ysQWVk7qUDldeYFdd1bDEb5TNL367iBWka0+gp32r7bjD3S3ieITb3gR/
WlkkycVpZ9UPj44hkWj2ICUrHyENDpQrNsPKn1XFqKE/ZzJQzTej+INa1ArKq31MjncPeS7zytWe
CKkaVtcSwl8ozo5WJrniqoByvHwYM29NYTd382kiI4QkT0Q47J+tHS5wwRiw7YXv0LsNp65yUMRt
Su9OUDg5sP/9yV/HAQRgZsLh4OM8T8mF6NBA5DtKCPfLruiSm8788j0Pgk7pQ3rzYRxIYN207Luv
f9BlrwGZKdR0zfDcJJaeAGrSoWSNup8W28qc60PaUMUtmOxLp9LbfG47fTL5Sl/Mpea55VH9NndM
lRvKRHbPCvCsC2Vo79SsDnlpvM78d/XKar2YeR417BbIB5cGI5kqZEeC5iJtLeL/TERqxn2+dpoF
aayVUI1/T+SYkuRVQpcH8a1FIg5MV/eTEcIe/PygILJIgG9nnbM4RPgm9KK8UQgp5HD3qG7/jxba
ND+BsiunWnpbrZYh6wdZ2FZfvqVo2C3Te3inuqaHU4lpKv+fxgKk1KNN+jQgjEGIcYzTUX+PxG+D
6zm5R+dUwDMxZZPnfWcUrfv9NS+iPyj3dyPnRW6RVENpo47ctDee5lBLQkdstEfsuyjkb1v+k+hL
BpRtKd2CoUKjRqe2lxKTbIurxrNUVQcnEoubTcOLg3zHw3sQmDsjGiQjEzJ3K1o+PmNbrULLQ2fT
nqItDJUjBTrPC8BoTRh924z19+WQqjS/ixVXWKHgvJ+G0oz2BD8lBFED8Vm3XY1fTC2pIaZllCz3
y1mXXpwGvOjdZ8x6geI6QUnH6CKVIOp0A9uUAB8onrwf1qygksT+Erla0+xf7ABreQvvXk6XrTqo
Tp97Dx7sfphTVxHcBPGfdQXO5BVpMHrwiD9dvL3tvcHBYJIdoiK5atfILq8iVb7hyoRGU78TwWmq
IliEmqIPU9bmYOEV7SGPXWgitxYQ1/3eRsYU2kjiyWGEaDgnQz/9fxY4ugehQXCX9JyqKkhLZ4e/
sRLX2GtohmCczISwAsMP1NmrQRPxwVTgycTOPXg6GxeiPXc2K/bdPWihCT9uR3Vz8MkoSf4c6Rah
KWxj0ppds3UnAc/ldOOEg5mCdsGlNn+QNeITCk1bEt+JecNN0PETrMyT1a3WHhpX2LXSlPAutQEZ
aFxPkbH6kP++58T8mhfK43hUmXcnCYz48o6Qpi90er0ibW4D+oAv6A7DhbdfWZBL9vPb7rBUkNDw
ndTuzu40W6BzL/AGVClzZYKfit+ncS6+dCXu+f5/lN27FCu1HiQrq5OGc8zoq5742lALFqfEdGo7
lDVwKk9gCdr/nqahJrJfNfQ76DIXXfPCcaeojPKGG7HArmrIl3MutX3+EAkXQVQpjdU8hLsg9Kbt
2HRW/14G634/6EdHjPxKJUBZQ/eEBWa0i7A4O0/zmv7j5ehnG+4eoVjPa5RN6m4EUz7ce0ZTRdKf
zIJwv9E5xU1TmvXB0XEVbQmzv7R1IvBK7qBL8phInZ1GeamBnQ15wv/ajTvl+vkSG6QA5X7IvWHk
p65nhsUF8q6uRmDar+nqv1ttFv0QJle1uKBbKAjwmWVz0XwZd/ds2unmsgr54oPOMptVvXXbCLyX
Fw7WQHU3KS6wA89+z+twxjvosVCMZFtXtgGc/yu8leawy839g4N7zbeib1u4DMHespUo/Pu958IQ
58TYGq390UbBzE5Gszvi8qQgdRY1dHrPf1OlEmiwaIbsRsKX1SoYME9bePhNzaDRwPv0WmmpA1y5
M8mHSBl9i6KKYAvSZ//susZ1EaTRLvnqJhbUsHID2r3dQqJThBYMWgHjATO6mgJVXgV/xJCRox5l
UCxdRogkCU0PDroK8HiMsrT3kr2/AQ+BvH4/1enV65xnDH62v2vVh138/uXOM0ko8RBAPzopqPb0
Y+iUE5/3sTEVOgionm3NBz0uNywuBobBVYFmE9XybGonMkStnliS/g2nG+u01x55XtlKuqbTIQDq
8lJoP7jp4pyrQyV51UBy/OO8FvStuSlP5HPzLMdCoaJYEmg2hGtKrc4bRuM6rqwvRz/541m2G883
f2bcDShX1pSxJhYeQ9l9d5yBTLZVLicID1N+TZN+j3zeVg0YubJussjgyCsoaeAkq0fYskZfhgYP
Jt2SyS2ksVpwCMolD2xZPWDeCmdjJkdVKUS4hIoMtOt4HB1u325P6lIDauSHAEIIs+vLImyz9Scl
/ArUVvRNtmpfi9iHXllCAYLzJgXgIkINw/gg1uNbLqwTMOg1mO+0al/WplumQlyCBlwMrGFm56Dd
zzVYs4qq9nVbWkcNJ6E7/8fZv6glaKZsxH1gIjfRvcp+d3m9HipBB78RSit6Mlj3JKeldoOHwIfT
5TWIUl7GJ8n51hwcfszt/+EpvdAu+GXB+2GNBalbqCJPd/UlnussX3D+FhW8Ezts5Vk/M9cgfu4B
ZJcIbzNKueAS0/MeAyEQHj05UFpuuTbY+73Ub3y7el3+zLsPPrByaKY/S6lUR/1yVp3DvOkl2MV3
LjXOtxzKYmNl3mSZk5ybiX5yw+tm3D48tdPESe9uM+77GzsK3apFjsKCfKj2fAH6PvnZmySR3D0T
Tg3q7uKFco8VEmogMmmEmLBBCl48FGxFUFN3UGCGo9bBR1K3REY6nxIZPXG8SAx3OvvDkVo2Oztp
VNjOTpa68XUsH+eQ3S55nh/sEVCaTNAgre0+DgG9+WpiilLL/bDNB2DUm9YVTHEWTBY6yIXhTyPB
GqKdgyw+0fBiZyvP7GuNnOXvgm+mU8FmMXAmRRuM+8auwoJc0Db/8gakLF45g9Am4uc6G9W3GRYw
JVKP8nw/ZkSZG58MhrqDc1vVfUbBIWHBRrAR6EYRzSX44LAXZlBdnE5K2rHZo9UV6ZlZLVyMOyjS
0VV1Ui7cQj2i7+6B7HAsEwX86S7FZRe25Hfq7YVWnEWBxNlPJFUjq47ujEUwQuZ0ZEArzSInQqMT
dQedny/NHZZsV8CAgMDix0KYplJVF7Ul9ladSVKHw/iEa1eBU5bbHv3KtlqkU8miVAtXxlpEaSzw
36yyv9ZZnCuzVu2LCaKgQlaCnJf/Y66X6EcqPz9F+Smi9HiX7vUCx9LGY081vu6rdMg5z+iCqqlX
iw5dz21aw/3sTSd3l1Ep+vMSnVKsfoMQtOXZMYTL/fsfUWohZCcd/0zfX145kG9ooqpBp8se4bjA
xnv+/Fddu2KM4rAG2s9WtaR1ovcTGbl8aUXYbFFjdZAX/RU6SH4M0qls78983Az4A3eQ2E5wEsVC
sBoneMrVNOWzQLnvdO3MM5nPo+1fGWhKcj5eGSUDD/NZESDA324AP6mQa2a6yh+qQfaHAh3C7qc5
xKZ3CM0FWXRt4st+DWGTs8hPOe8ZQfmC/OMRYV6/yRDrJsFUamZeqYUoXk8qzseZyhKU97ySe72N
QOc7aEvenrU9G7MR8bw7aHChLtlTV+2sDNDFpHsAmfIUJiIELIRZ20vMdRGznEDz0OZdfAj9u6pM
laXklvrEwSEGwDTIDXYxkbS4EYgUIjceb62POguqe6r+0Lrq7FiTlD3NoOu1Z+YzLkf82wb+Qer4
sD5wc/ta9vRZbmMIWRlUhZEnsvlJ0pkwjM8X7Kan7/3JVn3TLRIB7TMQh2fX6JU4ZGNiRCiCWood
Sb/fuvcBaBkyrBvh5xrhjI9A3DgkXykEdGOR5XEIdLZxwCGoqPCyoGUMkfFvgH4C9SOorNYq3P8v
0n6p4M4TouBgjFWWgwZy6DcneWshtEpA8nnTeoWPFSlcH+pE5z2Q1E+P2XRM8U5+c+BbYmD+/+MW
hvnwUG3rbjUKSwjFu3R2vBGmc6pBUy4LN+35IaNJ2sw7oj99Bf4hKik4rJufgNeNMG1O/qbJMH1r
27QaTvq3HRJBGFqr48lznFIAQTaAbX6+NQet1h9Zp8JDMHDLxpfX7wnShZFOJ0/jo1hd1o59e1qV
YjZ/mU4KqCh9++PatmuOZLGb7mzDRvoAvNlT9JgmmsHrJMDuN2Zq9dIEKR2lrGQPN/EF/TSDkQIw
xXvkeulCcZ1BHUXxPn3fMqIShtfxbG2hTbkxp3ZjSE0axl+xi6b6d8nRGLL1Iw8cr5+pe21MGahZ
Q4SKHc0n3/AHPAbJd1RrOCKvwpi1HBzYVCTtjtMN7RfZAD882uNh65Xa5++LxnHPYl7FjSb/v470
e7qNraV4GOAx0BjUZ0nOSiDFkKVg9R2/Xd4UEZvkEzgEM/V1NG7EsHqyq6Iw/eKLxoFAuolyCVBT
YgUybJowmWweUqfH0STUHV67Zzr0maJIgn8FvdOYvRPQZNwPUXNwhgFKurJMs4z4PZxUIS5jxoxO
rMdKtfRoUxQRRZKmWUckX9BS4ToV25SBfJNgo2NjuqYo8LZjdFm+EiIxidgQaq1sreSlbNIcJUC6
m5FH++Ee4qQYT2oxlnJrR+wcnuhljhHOzioJvqixsx5A0BVuraedVCNEBuHGlBvhBaEfLoLf1ONB
nDMMKo+ItBhej4fQayUY4x6KBd/IOuqNyXrYFsp8prLguBq0D3czEYNxihafWlsJkgW0amAr5Lhj
fb3xwcIQx4PkCFNiNUM2n6/j6u5T0Frl9DUsO6aEk179Ksz5fjj92/fPQxY664kVGOtKmEN3Wgj4
lKpQuhFxYY7c8HBHiCmA0YIMIk2w0ZKdwYMNyjysCywB+PUBcVxvIywlJUHkjw5LhA4anFdQwEhU
lAedph6uPG2O5d/V8FL5mrFlifv7g909XwmxglgPpq5ZjTTeIXQ1sEQwR5puRzu1odUCkMnr7+/M
NCUYO6KaLPOc4EZOg7a41DA+/Rv1UimS/nWzqzCF7Yk584UyW0rPYN5UoblwMEq7/CE1QVdk4p/4
UdN5ixvJjflLrkk+SXFav581ibr5m3yDrGG0pM7LXXHfwu6tzzdEgKb7QSdK+WixSM7t3o43RcAg
qXl5AG21lUWNcFl9yq0sfBYIRhM5+vU3qqatzZUGeaCcZBsSnob4WchmMUqmP6Qp+PIxEwBOYLrd
j9DgXx57itnrj50wnOkNRTv11CEf71XwRgrzJ6nwoebLG34jtdAnbR8TdmgG5nX1U+EbL/+qY8KV
YyiLZlcFN4wTtNWQmgvjpT4BykaOkLDDVwZSnzswaslzfeHjg6AmzommfwAqW6ZmYkELSEWvU8/Q
VHUVv/4Cd+AneOZYij3t+TP82qqUGWKxc7+xL6Pr+mj21TFi2OHlt+9csmLp/KHPiG01Y8jJ6E+9
b8keetTnfSnyW2KysIr5BnECTB3Hn+mo+6o1mX+EGH3DIp9rcDtHYf+eM9PMW1KcRIDZRcSMYndq
cf6o+1wLlM51qgkUztQSt0Jabw0AUqQWuZIOaGAD9jZPuy2RUo8CzFHJ+8TIZz5Mv06EGpGca14F
NiDzEBhJ4dlvySRxN4rGPuYcOLmgTlxO/Npid7HSdRDP6O2suaoIBIBNrt/Po4TrZGcTbaoLWBMU
0FUe81LhNDs5vQzyOiFnd3nkgCl3eshT/heDcH5mlXxZFpdipPM0wm7VfbxSh6FGrw6fCPWQWo3O
R7UZ0nHo0rveK0TlR87H5Elr69y4dWFD2riFCQrNhuPEon9xjA0WTWpgnkT1Q56721S/NpFx1qqy
QLYex/K7Lw8cx+vsJfeGGeX6NbLQy7/D2eU+Dfk2/99YxbkxlwKQLrwiV8t6X3pZcU0PKY3B6rlU
lYT+sMjjQP1tbyNCSQHMPuuC5SgFj/X6R3zHzYuqNvI5TAnAkFTveP+0bWizf3dd0fpaZRngx4dc
ASOeD93M1dtVgAkiYZLcKzXT7Y/8Jc8qdwKrbqSfUEPsM2LXKJNSuau5Q5MhvISqCpToUNfkAFd5
eAi/WMd03pktil1qouB9QBfiUwGE8OAvd6myWEmgf9zg8LB969CpBFMHyjFgeuoAzq0bWHXtE/TK
jU53UdlYUlMPEtdQ5IfReQ0EYIz0JEKJywP6irUqOzcxrPsHjCnIliqPkK7xwNzKr/pbvTSwgJzQ
ceeSCjuLfQczd52h+mdv2VF6nLpz/HAIMCTEjzynX26H1BAnfHSuOh2vemkLh9b33J0D+zbBmrj0
exk1ZKuO4ZnsuKc5e27N8t2oFUyW1zWBZ6RhdiNsic96bYr89KMitT9n73SO/g5W9LXtwjckYqLa
4art4fPnNWcgWpOpV2A58yeZjYPKfQEu+DcAXU9zOet9QtafQXp0dgcJmAYxVH0EDSUtVgkkrxoQ
vyyPBWhU7I0+NnM6vO34XPbmVUo+tJJ3e7tAJ457M1dBorlTJag5UP8SAQdnF9jru+dw2zNm2LxS
ud8yipU8MxnEMMxhD7cZHbHPZxV6nNvU6CAN+VlfsJddXDbtZHlAehPpaR34sTzBPuzvdsELEmre
hPuQjPY5r092HnqdM0tH7pvbbhN5Rxvqw+7PrscIFttJXncKzIQJ9t7UKchi6ad0/OGRaG3n4sPA
5EdaJtqjgRrnJqDdehfBOL/0iuTEBi9EQzi6IDnxBpeR46c0XlLHoMH1YCVabRB694gomV7hblNk
hCO1WJIdLdtIkAYpJhi/VH1YSQ9NvPZln1TCUgrxYFg7np0Gp18XeMMl63donXQ2Qu1FXDkfA/92
nig5cQqZkuiVePI+47LjL/mPerddWknSu7kdbHd18VDdQ1dqVgzplnTrUMOzVn6eHk1zwU5+XqxK
5yNGn5D92HaWZDwbgd8UCqo9ep2RiREIAW7EYUX7tdUNStUxBwAWcXEdSFMnFvt2YQYuh/XKU0UJ
TbzbtzMT7CTnskIYxbPoCYPp6sVJgFDs2e+FbjLxkAzFJYWb+G9nKFqaWoytQawR6UxdWL5Fx5nc
a6o8UoDOuQ/sEYRYCg86tnHu/K46kP3s+limj+A+PCXqo44qBw3PxsZgIEho4nhU8jfLQU9efkJk
unYSkQSDc0pX6xDsl8zBiu+H5w+4t5I8XMF6A5rrc3ps9LBqUm0hILY0Yl3cN7d/k8dwO4GpchCa
YI2VT2A8hvTNePD6obe+Z1NTdVLXuy7vzP3K2gWh1ZEmzjahj5Am1Q/zmIKIm+wMB1rultduSib7
fxbMcz62nDRarkElGgs+70/vUCy3mj7+iDay/eAw+3ini/lMEfS7pTpCHsCciqYrD5OQJ3OYSb/z
pqtwB5erwPswbeSZDuUcrgYJLzgtOk6bgEyy2rzGqjqYhmA1Ti4dMdQHMAReoVfxK+/6Yyx+2AHd
pbNZ4WQGpHf+GXxZ/YVZ/Jmuc9cmdWbMquiPLrthFIeXppcslyHu+GdohMEdDdumyK2D5avk+XJE
4vUeeCuXBkWM3umLxBi1memM7aFdSqzOREHsUVFIFvJATaJ9Jnr7Icx9FRC6bwzP22pEZ8fu/MzC
DwBTZT2ks3wPLPxhrBoAjuh0iZhtbd7urQJ2mC9DNuUovdyK7VGBMdEmVTEGyjHUSKfWL4+w2HPA
BqoaYJ0fmCsv6IYIFRTvylS1mpmypWpYnbaAJ5cRNSZ+4k8nwA6ia8kYRVwdsMhyXAlFm3+4hBw7
bXMFrOVONaBmY9+WikbClrW2m2TnhMKvCUjhM8N0Tlhotoi3sEhNwJck76RRjNONa9sYqs87kfCA
W0Q8glLsSHbgHTwp4959A1e3fLgTx+sJFSmX5S32HkwzTGBqg10MyhtTUbSixWhi/bZSN0MG/bnr
av77M71erbCbTm4uWaSSaa/Y4RjnTatmIgf5PmfXgWdj5pHw2ySncGyuO9+dQp2X6nZIDTcM7aB5
ZNurdDhSXMQjOKquhdxQwk15Dl7qTyNNFmcVZwirq/Kq2rg5yZA/rbwiROYkxpIh9A1JtHStLybI
NfbzWvCoP4oOsd7fBHfN4dka4rueZ7HDIYHm51HIDzKfBYlmXuS0dxrdgEyJoIUWM9AY4AMML01y
qTScjp4X2WRNglI1AG3MPnxGNWlcK5RfkiiZMnOBxsil70lUgEzcGz8ZJYj0/Kay6YkO9i/RYE46
me6oJVaNRcmElikHk5WH/Uf2+2RjHePsmWqlUbeqTp20UpXPydA2E1hPuJ5/vw60Z3Kw7N2em1PC
RPd5P7NBPb5E6BVK7kjrQ2iV5Qi/HpZCDBY23BmCpRfcJ25ZtIvwX+upc3RcWo0BIp6hWiFt/+RF
fo6p+uUmygrUmhxzhIExTf/4opzf4AdGF1MtzYlwELFuw0NxycVMiJ1BcK5eVE6r8uJ2uZ0FNvBS
xKpaBnxKqQRJwIFjwlwAMNUGVe66k3BvZz9hPbgu1kOECvb1zZbN5c+hTHriTOluZIjow5mAhI63
7WvHa4CfQxfEjFtDXRjOj3w7MfLxNs4LMcJbLeyHDvJ7Y9uWMs2+kzpnOx0reTfuHzwPKgc3FkLL
KPB6+gCZgxEsqW2BlKry+Tq/8etlj/UlZFjDO5H/3RuZcrieZ9hvdEmUFG7GRM7IL0BscQ/3tlx8
YBGKVjQ1P3RFPvd6szgh7kd6FVJHipkIPKWsUDmayib7XgEPCg8U/pJEbf2UafgznyX7S8pRq+RN
My9u27CqTSc4spPN2xNAuqrv4ecSSFvDUc6pvSnTR6s+BjkdArN39E+VAdEtO8hOlnPMrrl73MHt
sUw6mteVM7JMZJvJ+o50NM8+U9JGbr0AV9XfmgsA5phyTT/+DlZG6uL6vimAabDPbtcUdmTcAyI/
uox2racxkhUmIam8Z5/8C90ogpuKatoApiD4npGcZhuZyfmmGAsR9iL4ujH0y8XOx4um1EA0rmtR
EntqFemHRtFNEKUUZhjSzs5cGq+KsTcEKCWttcOXmxSyWdOupx9YXJ/he+J5sS1LtTJ8qpAf4myJ
H5kKyw2474Ek6uprqe1F0jfHGYM8smJmjHsSmzjvwwuqMrK33DRh83VdxtVNs+jmCsf1o1XqLj8D
G/w88CzJHfrp5n6ZN1Q0tG3ESkwPLJckO9hF8rp9pkhsY2AQMK/hchN76Yhnu3WFKaM9tuZws4KM
G2sVN5ZVv8N+OppBgCUUVb967Y/JDa+C7v8+SXxB7TSpBoHc/qS4U71PN908X6qUyFjvlj7C4/xN
pNU8UxsSg2XC4kULo0XFk1YReolfAlApzauP6hpwhbtwNrTGsaKb4hSc3aUR/VpGY9CUXq6VIPPE
HhIUFE1n+2jvt19lx/0UAw8qYALvcybkR2BjpimfOFX463XthDNxPp0nGo74MlCAcEVP3tvJpE5Z
ZzUJe8Esz46LeRwASeUEu3nHuCHrV1PTCKMXlenu90ACUrAbb2xTqjMHq+w3jtzxvQXClrMNeTvH
VqGQe/tBwuB5kNgvxU28QK48J/74uQccQ7/qkrHia5qL/cYeMEfPCvJAXPzezywT4f/H0SGoL6iR
xb+/jf1EQ7cH3xHDRaPokKFTB4GSdFELo2CnYWYlzixH6OHkcr1bWAso2OgojqA/6ew9ir1v+kfu
AkXxBiX0N/VrpKQVbwayNYgCFFv4BJoj3bGLD9qR5GoDFvxJmOnG/JXlrl1d+OiXBywdPYzms+sM
MgvpXO1fIJWhH73ZwYP1gGYCYaIR9dS7RLTfBRQ0DCVzn9z6P2AsqiM8KXJ/NX7rnkQmCQ1EEncb
zuH4lyAc7cW0SdIoBPNQGl3+8EPhj3NeyyR1sav9zGhyqIZIdsumcsBFNf1GiRJDsXFW1ZF45XyT
K+31XwmLJlPhDH0jNvlcyT8Zeqj3KdJgEcLzOMNINAgjQL1YREmcTq8GvorvEpIX0M41RQ8Er+ZN
Bp74LrrS7BYPGamHVRPTultO9r5OsUtXWsDyKsJuZdf5YCOIi0v+SsnGPcSi/RFyzVpIWxUBxZ6M
CLFtwYd4LOU7AHVmzvbmX4IShZJdH5qKdwC6Qah3RCBhQxXgs/DA1K3yMhLV2OYvVaZpUYKqT4Rp
rC19bQ+d99UOKzG44WTJYCOZblahndLGFrs0tQ43+QoFb+vwVy+dM5uFfGiAzjRLphtG4aFfEf17
cZtsH8uZ/giQEOOzhgil+rxvmiEret/TWfVh1LABWGSc8D93ToaYGpNpfM+5sKc/thhfX6T9FSmj
d6eDio2V4hL1j/9HiMQSAim9f8eiQpeOjT21YKADnn7Z58ANLTONcTtfa6CuxtPY5rAbdbk6qZQV
Q8v5KpK+ejbRIVNwH6maSwgeYphyFwlJNxzJuz+/zlj6+j685CM3hEYKcl5SDvDUqh5iMiNXsOM9
XWy6ZneKC3uAOyffgm7wJ0L5+oVzzoORgqhjWzzBR25bu/bS9yse4quHUhT81HyHvWt3E2PPWOdu
T/VWolDK5/Y31+E4NbuBmX9My+aKN1ebUakAzyk7dH/hBEEHkpnSSwZx2lhYXw3ckw5iElgMqOxs
NAZtj6mDp9R7hmmf/RE19yyZox3G5TZ5CXAmw4l58166WPnzV6xVbGXaS/JVza4QJoG39wqWWtSI
WzTp12moDp+I/kbY80mDcYaKmMY0mOTD9y9fczw59DsVEewyolqDuyInz0a2HB7Jt/WpVhJoro2I
iPHAVcCZRsADJnOaXV2hyRMbLW8s0Y3dMrxAAuld38uVrMqA5CVGV47GUgAyZl6eMQJtBdslYw69
z5NWZDYMoAD9/cmgDmz3xd+YSVuk1/0b9oGfOdjMM8rFiEyvvIfiSUwdPNks2yOrXjLWHEPHOC0j
Fp+2pegm5ybYDb2IM6WF1Z0b6se2WUd+NsIASm2oStkipzBDtIfGLDFS6qJd7qr7aXPQqf/Nos2j
vb9Fe4gIl1TubvHiJQHbzzmX2DtEI37u/8ckiEN6xjaF+ocfmsKuINsg1/i5V1Ryyr3+SoUtuysD
YYqe9EdmakNZ84ffSsbhBanwhBLWNo3HGiDbIQ6ury7+mdaVnhj2GQF8fxBfxpbyphTXM7jpX7mo
dUZsJnX9aas19nCfS5OAru/v3/dJCRu7/K5Im4ciS8w39xQ2a7qh3gwi8RyEaJE/5rTgc9BSvKPQ
77H1cu6ih6s7i0Kt24Q5ynuZwh+L1SCmrzK0I45UR2EvpwlLl/YflEaT8EWxvTdmsCZ/HXsnGo6V
go7e04h7C/tjDKukt6bIyAsFX4vORd/YI82dWHaTc4qY6LakUaXJu557l7MmkGTRfC+L6/zaex+F
VwVo6402OA/G0TjfPmuofxhICMYPIJYzmU9cSY/W92Fsth1TWOkZCsKCPf8obEEp01gkThI8MdQf
F7MQ6Cjf4FkqylrIz0NIn26ccqsem9AaT4Vakw8cNFQ6bbMp41T0biDMf4nAlw/qbtDM6LGYKj52
+nEVPoJHUzzSRZIi/DMwiSOhIMrTWcK7Dv/0Fm0bmaLLdeT+VkXvJ40Wp1wkN3kew6tqCMvg3g1H
NjHoH0pni5b6EiOrQdma2KT+TgRuMTU3QGvNyvCIRJqhe4CjpmaU0vF0ZzBMeZiYAQ3vrfnGxlNp
eaazoY0ufirAcLogPZNnf/Yuh+jBcQJOwZ57xKT5TK58yXBgWVc47O8qGeXkFTlyC0udxPoUTvMc
uT5eb1grbbL7gQxblI2SYDlsTJ+2mbzkd75ZGw3rqfqIZaDFefoB+r/5W5AYc78Avs4UJXQgB2yB
Q8feMvFDdOjjzrGqABR7MWpv/JsBlVqyCrjF3xVe08vzLZGfwA/PY1CC8TDYoY5GLrtH7/7JDQju
3PZ0MDLnUnzfCiAah5xH2Kxj3BTtM/wql+JD28fTRQkoFgWPwgMKM0Rxs+1ujX3izjvge+nKXO+y
KEpslAaeP9SK6XGJUjWrHRJOYTg6fyAS/MFH1KdSJ+reSf+KEq/OIdIf5OtBmGFpZXGwXm2Y73T7
RJ2o/7eWET6YVk8i4ZtgnoWoAisyuW2RMP/btxTo5fM6nG98p0RTVMp2g9rz2LHFag6a5M6BHLcm
4m1hZi+JywAuz9po31YUdynk9NI1tE/Xe6WzcIS3olwwv47NqwVHBtay1jzu7YVI+oo/XilN7BpD
H7lcZvktaDXi5B7hz7Zn7UsZJI5nO+qOLbyXn1pTCjdqxZUmQK1jVhwCLgDmEe1e8BTXMcCmwNOM
uAEpXMUsUxTTqcYgdXj5uvC0gyNWZnCb+gaVaWppe67v+c500NLLx4vzW3UMLXPRlNb63v8eD9Qn
PA8T+CpA3EnbfbllTfh5BG+y2bqfw9AvaOCsGEo2kJqik3Ef+jN2NU6g3X/z9buxpIqpqpjDmKyE
ptubxCxS0wiwTm4O+Mp4vNUVaQEGYRsaoIN1w7JulJzUeLVo5t/flAPGz3u6Cxo832BqwnPinBth
thWBkiYyz6PB++S6sSmdt+VHo8N0IDl7nmVPV3FAE00H1k/RXRW6JpvD0q2rH2I8uLh2czGSTyyx
rf+aBImMMmKLhPc5Hbq+WLW2dntVG8QDnFot4TdR2J7e4wEZT0IRKBpGQU8IFRkhVqTjrm6HHUiB
0sqr6v0FRC4q1xYZWQ1EDRGKStsZIEsHrObBnKShYILquStUAbdcjyY5ZyxzrVyjrLKVccVFTFbq
nNVNx0FgrxtduTjd0XK/VHQ4emg/i5eoWg6UCCZJ7g6uqwla908I/HTLnkkmov4HmDk4Bevujkff
2ubp0GKMatCPZC4uZknqHjYJ93o2EJvFB/nqIS2C8dwXWM0TRXuSv8kEHdFLeMFF+jnj3OyyBkst
c0a7JBQVdnZfry27WI8shwUQzP5de/a9AVgwbuFL/TqcOKZPGRWsVVlCzeDlxTddlZGStWura2Ev
ah0HJPJsdVUzVU80jXGNMucN5tp0uUihJ8iVdY7wQ6YyJOsbPZWvma6ELQnS7ZHc4Cm8/sWH49f+
Sg4/oyExSVUeOXQyBS6fbpNNJeVOyPYQX/4W/G5OCesWyJrXj97vqRDnRXwH/6cvJZEB5xIfaebX
ZgK375e07kvivn8e5MLz1TX++YP1G6CzEEyGCfymubEILr/KRhk0djos3OqgjYiG5LD4lbjGkBWg
5224eHUkNXpF9lFYLMzmCmB3v3AS2Ug9K18tKSTvKkl0CyETaE5+5mz22W5dRQZNWqFhxQQ1LVhs
7pwPwfNw9Dbym9ybtbAsn/3LRSr+YH5shJ6CP+vp1WguFvQ+HexacNLBMwqlfbqnINHlk+O/WM4I
LYnxRMAoq2eMgXd5/rq8A2+Z5bb3srn7h/a+zskpqU63xUClXgFtKdkoQR1YBcxtOnL3CqN1wpET
h6OmUEQ5zG/q3EnIfm3pdzvmtlaXpXTnQ1mdzjyzNz6gBCZgoWImqHsSIEETcTFuQW+XSK721reD
amJiCG7O4SOYD7eIdXEg2NusgqRhShb0QgJc34XIhOhZTAGOYiv+z7AxEukGXLMB/mMO3T2hStqd
r49/DUehl1cnMO93kygK3SxFVqdkZUX/tNUpII4Yk89Haf+hzqpwioE0+udsFysLqNAWCZzfleLr
jX5kiRhDJmA0jU7J3NJ+eUbYu4Ois7Cy+8aIoMm/AvHzr/pak/P0Rq2kGOg0Mw5p7qpgfPzwJUkC
ALy+1pFqik9yEjwJp0UJgsTyydKK7YnXpkHhDK95+V3Rn4zzEOwO8SaVzCFJ5LTPyz5lHDbZPKmt
hoJzCk9O7zLIALn7OGReiZmF5hAqxfoW4zHNouE65wPCPFvXi8hH/iZH3IcxOyCWJB9GK0QbMEKj
+OfzE91B9ar3jW3ocpH2QxK5hKGHDXuefpVKl0BnTHa/f7KV882eL3GPqJTDypWs3Z30unGNo1WZ
8sgQ8KaAbA87dEgIphuGW3thSB75N4XiOo07LMkMvR84XBo3hE6VO9EQlhzQepzl3SjeOyiREmIV
eKFdUMhgBaRzuc6vdPFToMzCTkCAT637YkK1KrzwgiVgXSHajfb8tzlmY9kQTIz0DLuFiBOLjjBV
4aNQMbhVEx0xFKN9FJ2uIKm7GBjT58eqobRJmJRPgJoTjDQmr0CLIqrLHl9FfRrRwKf3gEBPbSBc
JbhdjYoO+ffO6mzlwJY7I0C6CwDIgXfNOjNeeWxLanZpXfF4KQrRWLZolHrVnrY0ofWrLjGjjcSf
vxEuMtUlDwsjEA/R9BvHnzGkfH/Ivse2uVS3pnIrkpIG7bbpBMfP81aPzFaKMd8nYOa8nnUWE3yQ
Cl12jF5rq26waj0CEiycA/+RShTsOTHHGaUElQ7mA/WZN+fvV0rOCuExv2bobZk0y08FJQciyEiJ
iBowiuylVAh1UqUZv5ixhNWiSPnw4afFLf7GFzkvPoH88iY66oo9hGt+wc2UNtV6rjAl7azIJ868
/fCTyaPQo7PDX8w+8UBAivpz9rvieNsNvXuBiGIS3RlmmwHFEhTwa6cNYrYt9tsB19ZwPlTcbGfF
PcU9UB8NBBpFps2LJaSAC4MhSCYb1qxgHOJEcp4F7cAFCrIxWUUFJ0A7hDVgtHJqBPpXt8X9OM4w
u0EgtkaY8Jcem7IN7mj2X6dwqPz5H2GGv9WuuwyjwnPIq2x3P3ygu5o9VIh0UKOOeAR3OkH2ycfn
8DBWDnHmXCKlGKgNLCZNQvsRNmzXVncQVZ9s2RQfnrbV5ter45FZBa7f9JdSaENN6r0KwAePm4uy
Pr/KptfwrrMgm+mMfY+Kj+Gh/YUgSaEiHwbSSXMQJ/jdgOz+3Rj2T0vCcfySiyaqMl9Q8Z9Mxo07
mBJAN4CDFte18fegJ5VGMPk4G/SlMTclbJ4/3PYSW/Vazk77AI+KUBQ6RLNaCHzCy/Njd7DWLYEq
1SDir2kz1dlaZxFcFvvmkNjY/Dcxnq1qqw17/Admrv/PmjlGMe5nC2QOS6KJrpRDqeTYUlPHvsZY
y9QitfuY2V82GNK7nOPfgUC/yDWgHPGGRUYvpDx6oi2kuhgal6AXyN+glLljBTqhQ8W6E3zaz7uB
GqzvQMp1RvbczzAp7NrM3G4n+Krq9XeYAwj8noTtaKLa7fTqbiFKEIZzpW7j/hkwpw//z3/GhYRo
8WvMosgZb7tVh+jT9BM5NfgFDSF4b3ZL4nfUlIKaMxTlO8myzvVUVnLgys5O6H6nPJrIZP57f3LO
v2kxqB0Ny0TJi9RjgZadchSeo5YaAiBPJ32qOXAX1AGXh9FeXqyMbBXhs7sPCccahPxMnOx969T5
200P0ijBpckE5FmEPWDpjRfAOt5NBVAu/oUbmgOZDzBv5ztZhHVSZ7lGtH++5O4VwM7bvh4smprJ
Mz7ZTY9U7cdnQomsJn3gxlZmmMlccv2BgiCePer1YVB1q06jtJD9MyaZr4XpFotQCY/7qSJufQqz
uqQPyqGp9qkg1ro6MEEaJSQfQ8mElK5FTzNwQy6pc9d+tRb614Dn4FTcybnRzE1X0izh8rbcI1CV
BhCwLvrocpHGe/CoI9TCkF1NmzR4s10vEDchs7fUmuPvht9E5PQc7jDP+Aszo+sbnd1kwqWxJfKI
dfHvCQg89qkEIfDTlYNhldIMdynvWM+is21SZbsd5SiqpGLjUZYD0Kbi/xhYyu6wiMvVOo0DC0VR
GeQIsNR0+dAQ0rFDDLynkXgnyn16A2eoR4aHjUBUBOKaePTTU8JExbWYNj8BreMjcznZ02KlByfs
yxlHlL3ujJvAaiJh9blEa/Sbrkpoly0JjXwMdHK7fJ4NMNWLpqLeywiZW6nyR2mncrNLQDLYtaR1
7l34peM0Umwo6F88mCKC4TmsK8fY0G7Kub3p9JEH0RWgApcXCb+WFlANYFoRy0f3MdzsUOpdhRZT
QBDantq/bYpsF07Rgz8UXswXJk0GmI7vvSUerZtqWvXF770pFBrvYegsVQkOZyJq+jFog5lDVJWr
d9IyzHJriKykdnZ6u9ebQw+cYtOYISSStSr3fP2L4QxsREi1IR+OAMep0QZatJeQlU+MOvVwxt3S
zO82Pvt/6LIzpm9kDzd7hzBw6UiPR4f2wEpDPavpetWTMXNtYihqBo/nMBGUCXXb590eYhnjQAKS
Uko9JzcsHR62eXNOb2ygPfvisO9Rj6IvwS+GEcVfsEVjGeD0E0mna77voWQVjy5xnHVm2EkRa3Of
RxYk0zOXWwaxfl8OSLYVz2EMwRttmOpunIepVLfTNAAY9f4yCuyhPTmF8HNk/gcdJEWsE3UObAOE
SQj8HYFlggOEoeSzV621/G86pzyINgw83WKcAOzCi+aVoMOsYFobNhy5zZ8sHp17JqRLwuqKANfi
Hstm6h0lvl6R2q+VnezMXHo3Vv954wsPJbqKnxOYff0cp8G8qVgQ/KCfoLdRYyj5mIHzkv+llOYG
hE0H8b1ez+xWMS0zG+GGB5YfNSsORLpRsoTvFhN8VELTsGyoI1XeZWbndS5bfQkx4PCs0qt/e63M
ya1y6PHpAePBUvgqdZvnNXc/FqhCQPO2QBiSdmm71NsbMNTYM0KM69137OhIQcYGRCllNxKIJkHf
8qsxUNyx36JMSu7fcDXTQL3aWyLZ+/YcK6bgQA9Yw5rSBEEPvpjnmI9O1jHL0BHtp5Jp8/DTk24+
KPm4kqTwHz4ACd7BDPaY1vYytruU06oImsiB7/Iqd+eZL5bcGo+o0dE2VQ8RuKplk+rtK9GS4Jnl
e4SxPmN4jGiIdznpYhifk6hMXTQscT+eFt+SFtU5wz0hYe+zlPwkBVtqjCNRe7+KqqPmNkPMc7FX
brTbinkEJfS4jxBnjsjBrdYh2kjn1GrGZ4coU70g0bMUDdJZ9dWY6x3SUxutkdkBmwp4LP1PnVex
13evygB68dmF27EqGI89XwTFklWs2eRQUpPrliw9qjfWMJkVQWVimEvnJa/5Eg7uatSnb5EUT6mg
pdVnwZDM5EVHVxW/qQ+GVh7Nh3Li37qcf6ImUydqD/krqdQAvUC5rJ2yYFp5IP6ZhLOnAQghXFcd
c3sx86nTkBS96LQseQAX9AtP/AC6B4Cu11eycUIxIbjSUCZc20AKDMlsZTRx/pRLNyh5R3gvK9Mb
5sVX5htkPLC6/bJHTJh6CVIpT/MQrOblsYzZBnwoPKgeN1x2frpcDyAH4PsmzxzSOk6JjgnfSTBq
2evr2NH1V3+HBT1Gk3Ec2YI0uxcgDSOveHxsMbAbeJOeeelbdxe8UhCG2Jlk8VFk0r6BguZiFN7J
iipkV7KT3duqYbX5M2O9xYTQIFnvhC5oDPYaoTVtKyVxlXGF6uMurubLniTfPhBLHXL7vhvdHwoR
+6XS5diubCsQ6Os5cFA9DAqRz9AV9o5vCDSGYZ8abbgavdVXUQqJzLD2dX84rPbWloClB2NMGjiJ
+0kN0qZcq5xfNQzkBTWaxtUQjFiZZcVX+VeazOjSRb3jZzyvLekx38quPW3KhEFbo+awRbCAtGBh
PcWSWGfJOO3FGXCUPqWyIQr/bCi1c7GErwFynQ6NsUxunNrpoQ1uigpCzoJifPmqF7vCxsm2eESJ
22dAhREKoYg70OOAZkyh1mtojdSCyFs1e9qmcpq8ZZBSORXSTxcncM7RX3V/1Xh4HUOcfhf8Pafi
PeEffpbA0kDsdKiSXNCU+KJdL3ZJVT39pi2GXqog0whwfyRoB2CrC/nZdccgZ5Xfu1ZwKjm8yQ0M
AHulUBz/gJtJYQwbCxk9deb58eAHCBE0JGdyTM8bGBMWOun5boJLWNDQih+RXyT9Ewpg42wvjV6U
p7RPjbeMLCJX8y9hW2AqfVPPEGNW8Ao2V9NvKxCjTox6JURhGjoX/V+jxl+ItWWYWvaRWuPlwZ+r
4+H6BOC+8ZAA2cgD2LFIzoulvj7b9DBm4zlhW6kUgPQQUlINZ5Ir9GvD0EhBGdnpQkaI+aZuELhd
JzrgcQr+mXxD2InGl4A/ktbbFpi4WpDDqQnX0Z+kc/YJbauB2OZSMuc++hV40x+kXdJMrfezWyPc
m1K02iioEBTOc1jdavkbEo0hChS1oAKN81Avlf5o8ZpLVaiXn2eb9Ru46Jq16CCw3i0HWadnaL2k
PIIUQ5GGc/x49JAjE5JnKAHjblckox9IaL10dbNlnqoh4XQvGFSDiMxeLEhWDujO04v/vRX7crDQ
7sO+jiIptNmDq0BBQCmgA9UBZN0AWm7TOiMbN+8fzzwMRMkiVf0EuvgLF7F16qm7BVAPLx3wYSOq
9OEnmlz210t+FllF6BjKbPPkVRShFgSAKM6WwIHpxlT3p2iOk9Syd1QaA8rRkwV2xkUMcROUdXAW
+XetMbi/HMIFoBO3quezH6ebVHzBeWx5YzEEKCzpYT5zfHYJF6CPusVLaPW5VQFVpwMbZwBzZ5jp
Q6d6KIQOoz9QI/sBHv/uBnWkIp05Zrxq7eNmY22M24NiPOmEEA4lSFDLdtiq4s3yHzpt72Ltt2gu
pHzS5nO8sQq2EYzKPBGfcPY6sEZnhQPGOg3seTDL5T9N3BTQlKJmdOIpe7F2JUmh9q1OL1f5Eh7w
PpC52YLDl5ZIRal3yq4Pb6XUSj+4Dep2HYRqbJGFdwaSxXkqitUGxGXzxoh2dyoUppO1QawEJElW
w1JuF2o31L4qShjoQZPxTS2sD6cT7VxML+/5rfqvX+HO2QEgQdPphbdFcSzyZOevPHObnvEW9Qvt
YZYh33b6BaBl8LLnKQNFkVgBUzlpbEnUbtvIMpWqR7K3pcNZI7Y1LqxHDb6IBFMhLc7jjsAVO3fc
xwePWMv9ae2GAYVwgasLo+qc4QVT2emKqvscWhwCkPR0/IM/whKzYU73cmlgJTmE1pzyitXiVxax
g5ssu+CcyZFWM8pbWfjJUaxxHTJJWI58fFajg4nDuoq2DSYUhgL03nL9pZqDns07504lo+NZhRZT
UjCeczTtVU76Hn5xDqTWYQ4NsjfCOnvdfBdG/XZiY0HmmeNpw0zZT7dxZ18TURKwP1sQIeMvckei
AScfslFL8dNQrjyUOqAGZXTwkVOtulplZwD//jPiJA0Lb+uOcRIFKM2FfGkKTwiSKabuuWoHBWyY
PidOvcdrXa6FQ8chev400MblwNvaS5/MkRGu+MFPpNJpoishuLXr80P7w7X8D0imkRpSnOfrZWKl
3LJe5spkZv8T648PorxNohxLTh22u1S3w0hPCXxKa0rrOAvZrbj0aiWamQOpUqwv4oQl6FXvQBZs
TbYDA7K0ZlhWGffBMSY9hX/WrSBbG0iNiuUobKO66OLHQ55i/LRqNAcgJGAvZKqY8M59DWlgDSX3
trDnViHEhTdpWkBAGJa7S62h0PpZgR6bFrZ83XG5sSLHhpLpw7WYGayhWL4ZojJdH5+cgHRIxgzV
PY2RIUOpwa3tuwTGKUbW0YJUyXVgnludzcinZQxmkvjtDcLSfPoz8Lx3CHh1+5h1rvpOx461+w2b
St2iNV8Bt54U0x6xYj1COHp2UKDN16ttOvGYuPzk56OE7a55/8uDaMcvcm6yX6xkkvrg9ghu1UfL
IwbxEJQcNtzkEY5GVPifdFfROixOoX0j64bzNkPA2lI6vsrWcqCPlyQEgrsaD6dHL9rjzzFTw2zn
iVgBr1P/cW0qCwqnLOBgeafJogO/jbqFJClESwZpcVnJw/njbQXmOVZW0EiykEkcc1BLInndohJV
QxTZPldaYoxW/IueNbLUz1oOZo5t673awQ8XS0eKdoJt3c08db230hlywg/mI/rQgvnsyLi1G+rl
etxHjeBuQcLFQVMbul3e+nvv1I9N5bFtO3uOwYCn6KpBauW26sKsZscDg4SkITE9enlG6VBPeAEF
8oVXUVEQJlIEEuy8gfdmsNEtcGGCy8qfGCK0N5gtYAnZfFwkoXUaZ62bWp+VeGyg+XvADhgZEs9P
ZQtoPAYb2QfMLCtPrX2BxXde/ulADtXVnMtMrcIeFnHykVhpV+2cqWoIBJPpfewUw/mU6Ux1zS0V
7qPhipwwS2O4K0NXNcD0vrB0sP9125gnSA4e/1b695dABOF4MwGx9HCj1/WI0GcNEJs1v0WLCqgK
jDq2StOYhRm2v09kRD/My1E1gJYxDR3alTXCMiZk55c8r2dzzunEv3anUIdif9jjkvgZtqqpxI7H
VEgbP6ZCfft8t+r8AC8J2oA8CzV0COjpDHJ1+rTygRjk+zP3mhy9qI/2VmwjbHvPqUs/rvNjPb7m
XqKiDQeHagmuhPsZ+8FqLN6fUL0qW1OTvLeeDKe+KoBbg61BNaxFiWEuIm4TIeVDfi4AyPcpZmAJ
24oouqBdue5owXMTUdFUTIsPiuCxYNpYqDnS2EOl+51z/DCff5P+ur7GNxIPoje1ttTq2jKizf4I
euT4cRfjHJXSMXDt/Hyl2F4x+CJ56hmSXAaW1dNeSWtgLX7WiioH1XEdeOJkXPtntVZ6+2XlGUMl
Z2nZ3CUtjeATKerAGsu8mjK9TZLx9tKzdb0E/4kEoMPL2T5QmoAh84GFsf79cB12IRQcKUzIvgW7
WwjsqrvrA2y7Stv3rwDcwvYqV0s+7xpZtAU3ifLHxg0KdfH1ghdmShd6uHlNLMF2njKyb0n2Glar
iSPXiUbpxCGMu6OuS7x260w3D1cxdQxDiQQv2hHufA5ujDqKRVmc7jWkbshEce5ynGZrj4evVWDY
olC3tG+ZXQk2cnobcwhrctE8cmMGPKlmys8C+IRkSMSyhYcKzfzjbHRngPu/SLqzwRgI3zday0Z+
Mi38TzTqFpMB13rG7j89hjmcxP3r+R7NPOaTQHgwoCt2SzYuk2aSJgZTrPlUcb9m8/XuhKsegovn
RSyjbLcRCbe0W+c2348vN89MhuoKPs2yKwOdGcwcwnZ9NNFPpRX1hd/Icgxg9eEjqgJsCBZMLxgj
2rWHlHARoHDacJm7meN2v8Z1AK/b8noK/qRNRagq8gWxNYIu/Zw00hA5FhoAnG7H7MQ+tgImUsZP
GKwUPWskKecM33a5j97IiemcS7+EEmJzRj2ZgfGIvBnFaZP3lk9lpuQY+EGux7jK8rjBaULF5NvG
REryAm74jNylms7r5mYKkD7SIR/AjaVVLC8KW/gMz7fPOSVxM0HfIjOW7l+HjqWN59D6Z5810Sfa
K3CjHLSYKNl46hWlsohgDfXLGCe5yfV+qKenlNdWhh1A0hYtZupwS4swqHyESInzbSxMxmj/lMkb
9yVktGXn6Dmml/0IMyYgj2D2PP/OeYpSIwYeEA4rsXt8O1Yy4SvEqRR6XB18/uLaH7F6ahhFZSFi
Xes5CeYavjiW0SnCx3WaYoSVMgz+W+BtHCLce3EIvXImE8OXp62SusSAzUWmSXktNoSAauwTYJVb
xAZwQTetwHe7A4sQ4JmMz6xNAwWiZZ3wnzYZzxlQKMS8I1ROZEd698ctFOrFA1lDERZbUSn3VrgL
RJ8zTja6wwdQTb5E8SppFjKz+Yfw2FLWwbIs2D8CoOFaVa/JNvK8iec1bB+AqB6ic8NFVmf3PJTE
eSsrZKmztCfgyr384eiyZ90QAMozZ6DHYdQ7i3/UvYfbRd6n4kvfGtfmqBcO3VN2yHULaYW4RWpZ
wZK0i0kCXccheUNY0yPE7l082EiqvT1JTXVrjqxqYrrg1YXPic57wpXElJngI7BokZB1Q7pcAjJD
uGa+VwbNrJsiVrtOELW/FF5hZrspoEWT+fdIzQurH2A4DqKNHj1U4aKa98aPiEtWPBH8VNkngEWp
iGtO2avld7cmQlDw4GpElm0tvF3/PrG/FcmP9RxrzdyKHxOl+1t3ifN9kHEZKCBkZzX+4SezMtF5
Jcey5PoHiSApc/9M5LiNwbytaUhVcjLuTHGvdiFYnt9GCEH75JESg+l8NREB1jvY+DvHokiGNXfC
1fdrhE/tRo3liGVuwic1YoZNa6uFXByyxg0iO1LhPaaOAuOEpYA8IkaxxOhggofKQG2RXG1tswfg
37BF3osuE3KaeEBgreAZTQ1JO4TFzsdTrGQ+5gYVUtdnl12dcEEcTAGWNoKAcxhTABaa44qXsSsX
mAnfTCIev52ADq8M0z0DE+rgRwO88eVVOWkCCAFRzrizQnPrXCFOEDe1czgDHlPzFU4GLv59FBXG
P2l8fVj5NxtV5+7p8qc9/oGR8DvQjwCxgpzplrmDDxqblLRRt6ZkRg5kYKwYu5jqlLbX9zv5yVpz
PFpEAMSCznXzjQUgvml+ZDcWb2zb0U5Jw1M0mA2U088A7m64Cep6biRgSsbU5Hq+N8kk7n/5Bsx0
YVCltHXVt6y1FBCp73lVLBKNp2jrMm2s8RzSrd0MeTNdJ3OyRDHfU4YrSjZfY0k+ZQSE75wuzBz5
RnhqFWSWlTt0vlkzmEpsnNvTcrzhAcdx1LW7aU7Fgliow3ok9aUqgspJ0+Y3FiH3TrG1RJLXakjW
ICXBuwQQmaUQ2VkAMlraUAr/Msonz2pqUW4l+LGlJf2KmGJf+hspJygNz43/K3RZCugvqPx4gxou
pZbpCLK2TkCSP+YCPjBzdUaz57qfETFDAFXKwqAyIvP619uj+6NmCVxgYVvwO/FplHYI4fF8LvLl
M0irD+ISwpeqtJJjmiUuACJBRM5lhsspcpiyK9DjKhwEPEHhkRZToVtQE/5ruuHkVvPyeHYcxij0
+5ZYD5G1Ef0Ue3QM+PRPgew42FJVVKGvck0matFuu9ppUmKx4qFc6jhKbXB58njeHZarx7FcXxK5
eG/NmMsnY6oFrvELcsz5+V/R0YjGO2PDkOjbyA+Dx2VsbdnOIeV6rqtl2orL2P98p+0HA27AdUc5
T+/Ztp7J4+PpNlAedB0qRanYjHMYIY9cCQBm297v3YQ3FRazkBJDk2PE/8/+VgLEdi8aow4Dov7x
Vc7EcNA3FJ8urLCZ3Hu/VB4VuDptMQm04Xk5QbHW/xAj/kWO3v29AaP2fz6pKaQlI24xFMLz1Lar
LrlYH6rdzagHA05dhu2vYQ+zR3Gy2RsxUOmy6WKHNxxCMApFgrZFzVpYl5QoZ24wg1IRhEIXrC72
Dc9xPOsHZmqTVGiFAZpksMwgb+cI0ZYnuQn8TgfhjcACLx8CGumiU58fHZiwq55emgWtTxvI1JHm
TU/4nMn6LJtvQcWqZQFU66l+qhiHPS3MlqfuK2ZX3fmLvOuqJUnWeLuhX9KLSZAmtP1+pvfMvaCK
GpDeKjn2woReIN111aORHW+uLmzr2Lsk5Y+D9Q5kkaogKJCqf3xGfjVxQN+Tw8/rD5vj9akgD63s
i3osN5mKnwiXDTeCELTSRzPAODxmQxVza/Mh5BlHUZvvYb8/+VtjUaCt00KGqVs/OQ9tOBlC0wEW
ANZwkP1SwrI/NqK53uVvYXfXzIrD4l3Z3poPFrzUHeBBmdxHCFDwmvXRfuxk9pBS1uStszBY19Re
vffI1MIh/nSUJEfBw6T6asr1zxsrP14Gl/45Vr7WNuNjf+nYkURfCh5XKd0PYC/RvZ+aAS/8i2Al
I2orP3MBvuokB/QKvGcP7ENDGEgh4ZHldLnfCvI26EwlC5r4cc4aUI3ExcXvMgVgfacGmasbQt1H
utjKCRSavYNDWYy1/9vPkAVaISPDw/vy/1jg/wy3o4M93mc3/uDuVVVNrmLq/I85zaVapNUvLROI
hRScWW9s4wjGRS5hMXrAr9DXqjQ7cjc7Uo2u1BRjh4c2UCmPM5PW5q/hrNySoH2HRUJ9rxu6jN5y
nOmP02L2k/VoEThxqlRdtq7YrRal23PJwYNhcfYUGS9YpFoLzBwkQPqBgTBMeggWGic9fl00hNaF
Mp/EFUTcRuqUBLP5sDIPuhbX8xfflRRKgoF9hRSu7wrPMrYgEvTDgtG7cf4rAEGlW4t/xGhOkvYy
kz+FZB6d0OUCnkV55GQDSkeeTNvAHTZhm3vHsxVXqoDMXVL2W6sr92EyxMFq3gyJWXnVMVOnfYLU
itSLhgbQIZkPCgd9X+c15RizoYEv1+3q68BgqAHAjD2b+Ba8u93PcwCxiPJzJqcAWc/TcBzzm0FH
/9t8yAKvHgmsXmPGVSd6pVjRSWU0HcAuaT9yXbX93oiv+Ic63Kg8kepUpoVKpoaYbDAPH8bnmHKo
BFRY7KffTaleDlorLcEKkan43hJrzfKocbch3Pr1MkUXxAfUddKEtrBZ5qh8wk2Orq+30KmYmuiS
zcgR3Zp8K6uSIFSyuNWJcyTlCxW1bTjD0HQjRB8W0htJscoXaBSo0LIHxYBp12fLEY86khAsEJ8H
LGjw08eNkKsTDZZosFzHF4qs0v29EZuQex/VM2BD3/8XgO6ukBUPHBNXQgHNzRqJABPpDq8bRUd3
nuugv/Jt/ToOI11OOo+Vrxj2DmJ4RveCUPreVK59r76r8SMkZ6yXENSr8gC5rO+k6pWo8RYRdPVw
LQjcscE1qKg0dqivAY99OPZBPUPgk9elgtTjTLEKnmN0/dhW3T3ohVPfPYzVcRop2mItx2l4nmLC
X7wHoeWx+zlTN++y3MlM5th79hXHQ/MOvQqTCyuhgsOLmJDv6VRyxMeBp1Jl541NkbkL3DhP+VmW
olTr8WVPZ6NvMBxnz9L/F/z4awgPB094kp7kn/1bx6GbHZfg2tnlkTsgbYOVak2JW6ZJRvj22Vj3
pGvvnaR+AmoemAt9oTK6/Xe8bRmluB10u5kNWOCi6f0OOoYdGhy8EDDx+lLQflMJb1GxiuqGuiOJ
pOqAq2b1A7OOVyI1yjXRrHuRGIkYWLSbpXBReAyPQKFm67+UID097ohRWf5D/j2KdOaYXA7It4Ew
AHoUb5/FrWsjaiUMkOsGiG0r6fucCCiqQ2QUk/Mo5dz5FO7NgGfkA8rmcOqsVs6kRoOBiWceK6Pt
03Na61sluXtNYTb5xa79KYeV/q3WIglDIJR8YU/Invtmx5qhu4HCuj8nDVCUJBNL2b4UnnChiJkV
UzUI06So8/UI11hRh9cSdKX81TnUSWvNlU95MmYtfY5fovCIUj0u8hZGIE7n+H+PzrsupmedoTzl
c3BVklGDjmla2IlBNWRQNEHCruKpWIUcpIxHx3H7Q6KszLbvoyUpFXkLlpGiYbUd/OWJ2cV5HkJJ
ZuFfYc5NESJ4HUcA5mv5fg5GsTWeZsX1d+uBzWlz/K5TrM/HCW3M4KKPn8ZgQUEZ1xUdkJGNqltT
VoHucvWEq6euVzyNvJTLbAZIsrGR0cis0OpRbUxbLc9wVZeDpXnzNnkLMSmZIkhO/JFCV00dm2xy
Ic4AN1G1H3piA4pTHlQFtKL/IsE1oewhs6HcmTm+ATVBLZ47V1BAh4WNfc3GD/qT3K1YO9hkoLbH
O7zDKAW2/LfUOsj0+ADSpxDMSQ4Fb8xPVde0n7An9zteEwASbItcteNmTveF3b4Fr6rNz2K+IY00
GEuxx9tVp6fZy6Rdgf7C1jZYcR8PeZpaavOdUeWR/6gmBlUjRt1cq18bgSw43I4wg8Dy8/Bh4Kpx
HR/jVdvijG+095IOEW68pKpa3Xw2zwQnEhLYeDw7BOgYRYltXKcFim1Iwmn67XQMA/CVBlxWRnCs
MItbfWlPXJSKUH1Hj20P5c5e/OwamMXMMUe4eaKoFtwfPe/wZ6RvERXdfxfWQzMpZW+VpODcHv20
LX3B+ajeY0PSB4wpJbyQQD9kHLOvrcGzdQ7Tk5sQPF8mv8xjjJOIMPDiME0MoCuBX0QvsVQz4kd1
M1WUkZ81cD98qqSupLcQdnHoZJUOQ8GYfb/xKxPthoJsZU0eNeLQ5X2F0Rsfkz7MCf00X6ksEh2G
WyId/K5+3x9aZlYHAnui3rDscJXAq+D1tptjsKraU7EQbCnWSnMkadjFiJNhoaGI9ERgXeMYwiXM
t7y2MnJPGElx+vcq5rl+D+7Rb2+P9Kg7qiFu80+d08Y2eZ//miVSYigj62HLTH4NlACDbxbzlnAp
fJhuQDhE8IW2XJ9qtWHL/gwYcu7Tkr/GrVtryvQN6a02KS/C0j28AlbAEcoVNJhWIrfycWSqMiXl
2yAXFEu2zcHn0ncEDZkwSW8Gy1/II3X4MqQpbExVl8sBLNGuJgRSVsiaRd7Gs0rSCdUjVABV23/G
zWPYsxAM5v6x+UrmEpSoxM5ecgSF0gko9fSv7Pv7KgevayLh+iq4IdVnGRaE5DbDLkoueO2TiML5
fI/8GS1vT2cURyv+LLBODVaSnJzpCRWsjGpM7UqHWygcWBIRFLa/6j6TMIGvq+j8FXQGT3Zyxqyv
1ohEi3IIpX4l279kRqEWDXVGOPNabI+GNJcI7YwrXGgYtFVZhJ3W3KySZjpfQ8olhtk5v2Vn5tlP
ePjMGa1KRUC4QIHbEEkRJUkwuhl1Y5tiW45IYx4rxS45JbkAnFhXGY3yIPvDNklqqRTLGpaTlove
BcBzVVhnLck0b8sKXuEXnFCDNQhuvVVpWM+YskZILQlYRaumA/Ht9EPVxolm9bBQrfCXuZRnUd3K
Ox8ylMgE+73Y9biIwLCZK98m5DlciUuWS6TGEcxaAqTl+hQnXoOD4PxN8mbDWoXG5kpNIHvt+7kx
Jd9/P+5bWC0bQpBwN282gsetsk8TY9wD4heAd8q1QJ8EZ6ICPl3DgXp7A92EoXs3UawfhW3PBcnC
i1E1QGFzFxFzdFPTBqxS/DBlZPQGXpMgXU49XcsZZphEpCNCXsYQjekyUBEXsjDTniysEniTZnOU
7W7Hhhr62x4+VEVXPl1cBLC4wweteGXYRB2YnuRCZvmdt+HMm8j4EeJTRT2QN+OryP9KeoCjrWgR
ReWofZtmWJW9+1VqEEEzgW7OsYxgELbUbCIBOnOwY4wzNHw6XAGvdIKg/7j2NJEA4pq9LZcazKFv
70YU/CCp6twQmaqqgm1pBLAG1IZ01hnmiuZCGAC0Nq5JUKKMpiVMjWZTFT8wIrXj/Pw+hQUYyM+F
xy78YdQaCCLO3KNfEC03ZHiUNNMe8iJpcFEi0bXXBRcwiCZwxiB4W8QBQu52LaCN1Qa/QzXZYz3j
Doq9fIM9YuYRkOrjIDjiR6Ss8uWQBz9ZQGr1gPABGPwwBQN8h2AwY9NnPLtHdxJtX77zqsBwgv3i
73jcDX1RK9c3XlAUL1WwtaqLFShfdGXUodPJkQvI0+R07hPIuAN4d8ye1+riizMM4aE710psXzNR
bpQ/wRIIbVhpBzNDapwG1Lh5aBBbUbR3ocOBtZK+yD95NuC+7yBNboayfenincx+EglEY4VKLlwF
NoN9eNJQVvvNKKBDDQWdxjWvgpvFRvqh5O1GKhhdGz3tJhcUXMRZ/gkgvc28f1m0YTOmducQfuv4
rP1uonouxib9EWK2+qMxruiB2uUAje+XR9Ce+Y2D/biOoCp9vlh/2of0RLnbl/oqJkYF03Rlu/wK
sfBiLrOCqPZXNvGGwawRIcnN75bVdwvwktbMksn4TEYXd3vSn+qQusd6SEDtcMbVwkkRZX+OnjDy
G6uaj0CuSqNVHwuzobPZoCoH0PNzG6r9mAQEdPJ4dytRIaWWAgTPpMg5yFsf9scMEgxZHB64qtgi
npYc/8rqBDQUQM5en6LpaeuDxjWlHLKYQc/6CTLexcav1y/DXyIkEzTTQ9dP9NVPZC4Pzs6BaGaK
q9fTh+J4Y1fxLMYX8Jzsr11qTXDIWjLuCLw9mGWbhoQ7tfbz2drS+htxMKKlLATcLPxnac2Ppogo
MXx6nwCGIN8MH+qFhBfCEJZt01MB00FStCdEqqPrUrWm+08zCFLxhm1kOAeal+jvj9ycFpNqRX0Y
W7PUhG4+zohod+4iv2mJBovguJJsv1C+gOGlMp5Cd+ev0ATefmI0ctZmtdf9NZbr7gn804vcQNBx
7gGP53UZhnnpmyOy+eI2goRvrXXz+A93BGR7oTzY19E8SR5DpwAn5SV1Xzl17wwsye19YtnBFJsR
mJLmPHHBlctldkrCa8biHXl/KlB0hNs531gJgPg5DdHguTG8/9wI1lrFIdR1qvq6hPDbbG0Ui3FG
uwCd97gJFcjOHxAI04pYtbjfhP71HjVNphLGijIg9Pbgck1BIOOQOz0XYFdhQcfXy8lKrGWR1BDx
tVh55WrPIOMw3+UFggZ6P9T0EDpVrOLDZxK+iqgaCNlHLXni5CLgIvF/AJdSTFLJLAxvoq24tOcZ
w1JtMYGmWB6DFYJVnop+dEn4D1jYK1UK+G39QCP2ZRjAT5yS3Jpd0SApiZgQ5Xv9OmZK0RI+q3GJ
jiikmpB6fvwLfga7ufV0GStFSeW9JJUppHUs0Lsg4zcZdQoYOK2uHJkqn3Bi+VyAg997WK9Tleme
A2D9Ho50Axgb3JPNwPb48S/WqPz0LeyzjxjdIBOfsuKXsRYOaMJ0WLQjdIP6lAJbtTHOZBUb+Ic4
2Gm7Jptf8PrIv7Te2j/PA602eploRy7w5j8qN16pjYlvu3rXeRhigeul6El9OGtL8L2lJECtD7IL
efpmBYtMP9mAFU80eE36fg0bcgnLbXG1A80i6/OR3cWlJg4iyEXq8qCp/F6ezFSjUO1FRPVrW2MQ
nb5ID0W3Po01pssZQK8FAY2nUJPRBHTukFUEwxORoz5O2SBOwCMXKRyanrKSu+n6kBaKM3FjP5Oa
9Uj7GOSMM92ocA2TXTGFbWe7SLPXwltFJLADiCfGQStYzRV5LPvZaeYtcTJjnzkp3bpALeAaZTqo
poiDqpTxxxjgXW0CuWwAL4drX/r1qejPBQEgVSyKPCsZ+YDt7IsYCcf2EBogyJn52Eu/SRLJXupl
TbTLdfuRB+ZKvgspAIRX4icTOA5bbWPUOjhUPPdRLCZNV6Mz7M6U5+8PSKxnZ9wfok/zpMBT0sjM
rcfUCatVv6S5Z7TOorS2VoGYOZ0CxsqeYeupz46KrKUbA6XBQcyWmjJWCGKR/EIuxqaFwXv28K1K
cy3UL1WexGe/hb5EWPdB4nRjItszWUiX6YdiEiGxlZVrDEysVWvf6/OFXPDFiyHigJej3Rg5pj8O
yrP94kD4dyCWznNXP1yjgaHLooCY1jQHJqSqv1qZIUytf1qPoXqjT4YRsuubC6uLWnhPbFnwc6/u
PM8X3xncaCU4IIB0WOMfqgjcRhU8h28P0Mzv7EgD1ENzId0HQrzPDI6oNm/in3Hw5lwi3i5C3ill
1KodY/++SIyYoqZbRTyLEMGLtnstWqN+vcRpvs6YwMmVMHuobw99qNpDRywD41iVNckZO7BWIRAk
gusDadIJ7noBSv2sM1jIFSFbVpJMerIs98bN6GABQg04hxoJjyQ8w5G55SQRW2kOK9XkrAsHy4A1
NsKBzHPC6AlKA4ys+htq7pdCUyz9uJ5HU4uUiA4mW/O1iX4rTAmUDeLYek7MFeHVV1POHhfiU11E
XgqYUd2jI8EAUyEL91GWrIcJxVxEpPws7EfrwCP5r33vtAAsuSRET0cK2BRIw6kQZZDfisEtQlM8
7eQhCOno5jMcQyL1Aj2VCoXq8XQ1bdhLQToZOP1Y1p3COG+LKLNCGtfUOLZOCzpl8nTSJT27HPMX
ixs0XeglyOZoMFsCwChy2Z6uuG/YGx2RVg0OB6c8wwyGP/LtmYLVc9e2v+LpE4XZuuv62B3+2WzS
gEULECKbamIYw+B8aYCNPPBwuUoZ89kMGlAF5uZF5LDwg2lMq8iVE9NWTJRnMCqkgXSzGbBlVC2l
Ohual90WhT9symz6e/vi53D6+ylddvgy1xNeOEt+n8/mT+8whefyHA8HODTpPE9N4LdMdcshmDwc
s7jCtKotvk7kgAID794pdM+WJoS+tm7FzAT0NQbjNd6gLjKWtX+zGGVDMSYWmq+02qW/9qPnUUIj
SE0kE6NQU7Ka+DsZriC0uPMcgRZRrj+MQPRhDGrKcB1qFapx9ryrtb2+8ptGfZwD610bsrQrjBGa
n5IYuOeI0acxrnFQBpDsMpSR09HRYcMDE4efXmqhgZ2Jf4ia1c91Z73DqF8vrlYnPXKQKQe8/OgR
wMx8/AR9RaRQ+BdqiuacowMdYTOZNxKnN/1CDGUAUg7ecJYCnYcl0DzKExHnHvsaBOrcghCfPHd/
NFyqHOo8mItEYaT5PGpUhp90RNSD6RzGbakViC3ktNIH+u90bSot508KOaH9cVG1Rx12mT7rHWI1
uJ9WYu+Ww26E8uKhbFY2IFbIT1vrsYQ88lKCSAGwbfckd/LidPmT+953Ws1AlkQb/glbKp+htT+V
AhIDRyUl1YSneAVQUToRNCVaJTs/VsYkpyYFln/0oqhXKZO5/hu67ZaedQ76rOXFhQNG65v3Ft1o
hFJt+J5DGXcYLXPPnvSvJfffSNpe0IH+q/YagRhtK1LolVmZoONR/X6Hufo7efUOEKdfHngmfXYo
QulL6zw7PKbvL6zY1TXs6qRbH1VIFAmGfVHVKSnRNPsHIra0H4MLHyGJKY/3GxwxXfkW6PdE02sO
zCrsbGf5j+gKWTeCXEeEkB5zwuYYPLst95AV0hOLz/xD6vCi/zTU76DfNFQHeR4Efzjx/C0V90B/
sq3FNvbYzZbIF/mUxbmgCBTVrncQdSoXYvd3LUzYpmeZ+OD9KFAxzwzPhn5Ee6fEzggHpI8xahrg
Du4KPNVbR0zntILP8Ji2DvDhHLcMIZxEV8P1WQ4DlIwe8Doxu5L94tlo3SXSNkbmkKB8cfS3qfT8
tSQvFQ5jCfleWfulEAUGF46szgLuTCJNeUmTxVYw42BZhPhtIf8zYTPTDRl3hanzukQ7a8MywNab
ESvDeOxTwHHa+5pcv4lSW5wRRDy1ztgQJYTybUxO6x7bfmDCcmO1KkqTb4Plj7zi9yin493N8z9R
L5KizlGMobUIOOqDBnILoXK6Uyet+tJ3S8RnojfSh29p+hnLhcbJRESuHrNhCtzageYRlySCyg1L
ZHAZcWhTwxIKjWYGU2xPIXndvHP1zg2t6LyX4rKVYgGYOAOE0PUfMM5noHA1KR6FXIYValxbN6JL
5oxCnBNxnd9cEt6hyP+ONLVprfg5p563zNjFjRhMBPiMbf3al+te/ozODwpryy/HMdhr98akjiK6
24ezsXOHVxfTLU5X2nLQHfsHREBtmcW9ZOsumNUv4lA+U5MeJVLhwxPDVYRZP3rPIptxyi4bz2zB
36FztMKAdVAtqxyuQgBR2NaF6xdmGh836rqPtJx3y4EG7QltkNUD8ZLusQ1W0NnfkvlvuGQclymS
wI4pZak/ItmxaXs8NTQfrKnCjHgErciMu/l9+Bh3Yyw/rEEQL5tCbZ8f4xHilEQB842GJGvs5q6k
oj46MWqr+FvbWBVjUCD9Mtx0aDNOYj9RSqaG4XDGbu5FfVtwmKWP+V3tddTDPhpW+0wMbrH0TwUM
HnYU8Lzm+IJv3xf2Y46hP0As86EDbsB/ztlDHOWZzw0NAmj1KGCaFm7CiJnITGl2J4IHlr51c/w0
fQvFl8VIJWTnibUL2f7YOrRQhB4FFP2MZcY/rSm9cUwoLvdWMGs0lu2euOlDSNlXhsrNnqfWTD85
tRZclDmLB27OUShRNIihZ35lDFrRl3mwfYvHEd9pt5Xp8qYK5f/WtvEptlerdqA4z9FuiPpsErj8
6he4fz9ftGK/5d+OmvYKdq6MR/G6D+kXI2JW3f6c0QTFYeelLDaH+uf+pejWify0hOm2B5KKYGQy
zLSaWMzQ5UkcADOoyR8heXFszyULSMnLFibFulpiy6Y8o5tMEVTEc+iO/JqzTLX5zVDsfpBU7jjL
bZ5GsFTQTqNOojhEO7pV9oGpQYL3clfbIKkkwT6pZq6xirGBLZFWSpkbZdgw/h4vBkMwIjP0B/+p
D+z8TAxS+yZX4HVd2qvSUABon0SLa9PIxPv0gNGhBuggPVeeSam64NXebVnQ33kFHWeWTtSi2CAV
lpqsyC/Ygbwkp4FAqOxV9dF/RbIk5PHZsBvg2kcDI43CwlhVyPBTCR0ZzjJfW3k0D86ayMwv6Hks
jdgDi4CtNYkVSgieaG8vwicQmIyrTXjy/PMc74cSQy9O2r4R9cjqyJFuYZ+v6eLSX6iiLEGdMC3o
/D5LvXZVefIF7aMXVcRCVIQpgpsm2b/wOlzi4NeM0pwXhlvrCNuJghWoWbgTTuAD0+EGrm2nwhUX
T2H9Q7IySWAdeWJpjElXQ2QHL6UUymshw/tfiUQJd8Xg9w9WAq5EoXkeylTknzhe0J2x9+bjYWIg
9Nv6jJcovfDVox+94hxuHZTjucKjfK1wUkFJjLaaHaPFzZ89BHpIgZ3Fpb3bWrpbxnUkZixm68N1
9dms7WK4XQNQ961D2Wpx4gmzYz+GIlO8JCqJgrF6uQMisGsnUe5U0rD5dVexKPi/2loM3U3Yp9Gt
oCbJT9acYFVmGeSNJaXW+gRyRwwjbTWni6ZGTwY1vCwCfGDK0FKjpXcFlJWn0UCdTSuwJCoytfhL
9i8MAwI6H6BxrcUQO83Vs6wTtorVyE+7CvDBNi0xHrigDnuWIiOkzoIgBw+tsXaxhHZxIl7cOyQZ
z13eRKVlfpQ401/0JTHm1WoJRGkCKqHww2KoHtRidndX4QTkEa+IIu+B3oqyYy7wEDAEzIz6hy8A
h4gZPcZjszfTByS6cJ0TGYTdAH4EMmmNxLCtxf9m2pMyEsebUao/3ZEN8JqKxCJMbN1K/5qD0xlx
xHV4dhc5+EcdW1Q8pDWXrhB1s4493zUD/OrG839hNaTDktwanslgGneomM706g/FXF/ztUdcYmni
nLdRSiN8RYrGxjDbH4TUBA72UIPjbSkU67skyww2kLTgVI5vVoZ4h15tCcbIIwwWnznkCB+N9Mnb
PNsN0T5vQPKKLLrXNuGaKUI0/IwflX+jpvyIlBgObteAiJOygUv01oJ6Z4XB80hX/X8kNKFkOpwQ
NhJ/UdZ6tTgjRB7dJGTIEvLdubdPJdWg0qNaEHE5jBWU8flDeEgm8KDXFWrLtui3T6TJCUbx8DsJ
47iaRCSWaK6zo55mxvnF39BTAdhVpiUCcRaLNA9gIdLZN5w/r9PfJOYs0kdn7+4bk61Fp/KkZrB5
Deh4MUVZDNyJOk1VD5wCoP8LUEzEUJ0B0QR/2j7HnU28fafc3jkWY4dr42T9fv2DcNEfQCv4+8zX
FAlIrxONZBsNxPiO3NuVom3A1VEolIT9jno4tDjH9+qWYLvQfXkXb7LKeHI05Xu5vMUCq/0nw3s9
IrQxFtaYKiDuh2wn1fqe8kcWAzghsXSz1Tj38IuW/Rs8xdmIq0snt3cyVuW15xz2i9iKsw72AgnE
OZ6ACTJmztg4EknXowdFS3VsHnWK9o0D1tm825+9AWGWtL2mxMWR+eFeZzz7zEh/hzJIKRB4hkZm
QA8tj//qhOCRVKclgrmxj1e6+xCkrMWDyInCOZU6tu4j7uysMxjHl6d4fnFvvSDx/xPCki2t596l
eMN19AETOjDB5F1byHj4t6rNiuJomZNWRJT00dJUPhf4Yqwu5ysBPhyROtZm+sjEE0yFrp0peDhb
kFNVHkIiIUqUDeVWRIF0f5jQ0tZLPeSiVSlE/87b/D1sRWBKRwScLY+plEd5pH5/iDD3ti1yQsCR
bGtIeMjCHEBViwuWf6XQgg9IX4BcE/CxVIIRwKut4peqlAXGa5xybkv4Ivx5GJNceOBHHfZnCLrE
6sCqSQBEdd//vVIgUVw7GiexuB3Q7x5bK+Ri36EVDFsc+RJ+ssSEK9HDomGqtRi/SHQutJYYJJnG
gnV1Mj/7yuKJuQMLJiEM7pmIgJ1klvh4cq/HL5zg3Igr6tkUSY3gz/3l+vdiUl3KPwXURvK9NH10
3yRnNYgLk9LijWirrkVH2cFJDm+RD51ECYxr8ASwlI25vyYOFC6UHwQcWgPzoTzyUG1aAvDcHQkX
CXmzr2x54wqPZSLdAhPrU3gZY0/rfzHWvOJz0sABg7MMrrBevJeuOVjbvFOKgAfIMhuhAn7YhJMK
VuFCTy8sSmBxoNSGfqWtxD2oFDjhnMQg7j3Zrn35SDQH+xLtfGrx7xjKNiIiBgrZzsSjYp1xPBsF
b6JsxxnAsA4dfLP1tiKc+mw9XylLz2g/BSYG9A5esA7KSi2WeC4Hy0oSD1DRx5/kg+AecKdg0YOg
0vrAFjlOCo7lr4/C9qgQZf62y5H2TrfgN4prrfbmM7+070r74CsRRLEaPN1iGU8p8wEB+Muzt9+1
RJ2zj/LNJYxLyrwIpb5L3adxl15yusWa54UApDmXvuHOfOif3G7lfGqFMMx95ErVq/HVFLLFS+C3
9WaVlgGq7Kd9+12kPpCLy+Kq0wVOpoPSNHeZJtcUnFN5ibh+YR5xOrTfASxsdu67rVOUR341F4nd
htUe3Y1WtgorTRjpSmvmogmVScmNVMi4cOIm5L7QcEkpazalZRmnHjPQlKMf1jlnWUtMR15DV83E
zKvOLh+Vw8Mk1u5s0fenHDYo0xcj9JH740l14hBZAU+JkiE59EcWAVx7Cemi8n16hkm/tduDeOYb
VBsQnjlKszoWoWqncDmgN0k/vBPyzaynE+9yHdNoS/QKell+Kuq/SLKoEgraJuCkJG8Gb9yvyRXW
+H5XfE2OfTE+4cUYuwTPUu9a4A2WyPvqM6yT0YW2IkM59qkpeIISUA3nqgA9SY8+PXrOpJh2FY9c
GsCR+YHHTx9Jx6wqn6bfrStEWscv9SkptfrjshCeTbh54ZomwrliHBtq8oyb/4j9j6VFRfYwqw5G
NEJTPnSCrI8G3FEDBq1mAZfgBJPHobrFmOpUH2yNXEH/DqIxrevz5mAPSeHRtQIN0N+p8vH/qwpi
0BnXQnQh+NRtLrN6VJ01Dem8VVkG5UenxZATpZ2k6QGqxtnmIqfqcGdf6mq/wphk6eKEy8JsLzl6
SGexUKd6y3nunu2UrWWPiJ5NO5HUnTqaSDxla7QncJ9ATWaxT/+AJK/V9jx29bWvstNTSf0ri1TL
eNMYmxm/IPv8h7XY8BXVtpD2ANy57DcLPFho5kVTGRQi+dHm2imWfmY8KbPkoi+3g97IKZNt4Xvh
rgvti8IyvurE8N1CdFi1SxHjCYu4scVd6Mioy1GoppQjiahxcpSeP56RVP0hHLsk8aMl8iUc6/dp
XBExrtoIDpJNZCn9jiSNIMD855NssBdOgOyDVFUDezrA316JjhtfjJx5uJxPfueQ/sTjiyjUDEv6
ylzFA37XKxndgKi2z6A/jmp3hMAYg17MvFfmzMvNIlA9Cfz2P5tuTycRtqUQvlyXRBAvU0WABJ+G
bD8VpiUELaU8vqbYF7gQloCMLhL+GmfqfSDCKdAZUhLYEeRwc65ethr8AN09M9oYFt2kwiJa6qvF
NWdI5AUPc5xgTmjtaY/P7H+G05bFTsDVZQ8gH3B+9Wd6OO6UYQk8vMixQj64whvktE4ZZVu8c712
zfSZjN2s7RojpPDn/SdiZD1IX5p25yax76Gkwit/cG10xEBHcXJj5G9RgFKxpelbb6KXikHAfILd
zydqz6c7qOGc9ETBbBsJ0DvYULRnLJ/yUbYOjoUUVn3VmpBu6UH1bp3SnpvaG4uq9lGYw9O+zr+s
wKNY1wI2Nl8k0vdS5V9sb9gsVS7laI7j/9Fhn4pyqwkybtPLk2uvhmocNJ5IcVhIsMG18h2p9e/3
VqCiN6c5WnIf/yV8Um3tocVh2qKVqmFdsgeKZY2lsLovTvj7hZ9o7Xma5s0a/IH/i2GUg8rd4jtm
+QW5afsJeu4P9nol9bb6or+AXl5z+kMgDKmeIX/Z7IgWF/Kbwgt/0UVkkEhLpKPREf9bGGRp560a
GgcyYMragMIBfZjfZ1UL4xD/oOvLLsVqYH2Zy6YTc9oUKrDWXTKXODwRQNVc8F915laqT4uK2Lz+
9HHqVMOvOzuAjjo+x6DMcaLiPfTMkOV5kc6BZoooTREOjCCDYlAyU6zW9qR+0oOw7/H5REhNDwfI
yahsFGzy3ynwySy+V2HYfAI1UyX5BOdL3hJ2ignvBGvd0JsUrYW3Y+313nQaLkECNZ+qxUVLzASI
r+nAVKXwVvUXpImwu6mCHra2L+cpx4NwsicVnOQ6bGdWnVcHzuQ70udlDrlJBf6nwFZi37xcoqcn
4bjiCMY00PiKiqc5f+rVkcH2jF0OEXO6nKxlFomz8CpefxSypH6zF1TpD/dMcWYgpqB8sNLnIRzO
YkCv2IfTg7HFu0Mwidorl1t0G50FnHf47ZDeUi+bJ7ZU24f3ts96Sq0MJtX3R34/TfGz+YXtVjOK
3KMnDdNNNkDYmPA+zk3/7OmllHhVQvtxyb+1NwUTIo5w23pSpxw/HVj4Xt/WM1LEa0kaUA596j7g
X5o6/gHD2BfdDx7/54WjaNBilVj/GT+Aw4WGj3uixcM+XM01Ef3Hw711MXEQS+TiX60nVDDgswsr
fSebZBwTALXu/zomq6cGVQ5NKRPlYERepeJtXnQDIEKdVFjL8NFYIIBFFxgG+GorqccgdZ6OsW5X
LCbMt1WWQ4zPKPjxuIykVaDNkdzJa21wDjIebijGeHnRbsrehYNiHTkCE2EK4yoeq7XYJWA31Yrr
MaMisAop8DyOYIx/hamtecjyAuhHe7hs9O1r1VR14qFavTDeuP1zK3LhwGMgzW3iXD5red614mNc
Y1lO8ULYHnmuFA7qvQO4T1+K9f0PqaGh8W7Bda2m7NyWtqZvvrWXAXByiV/qhDe5Ltwqa3lF31XA
YW4ePc4KvdfV6geT74vmJ+dlZjYsYLicyHuGQjjIYoNm9B0TgX8ILSDwwuX1wRmnTcDvMVk4rADL
Twz+iDbGVbf+PWjwiMhlZQwULVAHvwWKiS6Ln7tyJkLrlupZnxYFxkGj9XZhZc8MgYz6nVN0S+ZH
e7Q3eJZIA/OC1H1H28cZOM/VlCzOJRhl9ubwYUfuX0KYXatYnhUOKibIQuzM0NJP2NCDIit4y1PK
qDGwM1G6NLZwTZZXWBNbXyrLWTBPVNpSG7Tc8ABv4Qyhfqts5zLDLa2uVO/AI50uEa647sbJ9XMc
N+yN67guVMv/TMfwjE4NYrjDVYdbSV0zG3ejrmDqIB1U6ZGlLMiKP91iSs2V5tPPwE+L6iH9o6rF
aY13i0W3DLdgG9ZzlNdrJaNJxkAwY6LWvZDC9nOltEITlTtCYpS/wxPyNh7CpkWq27e7wkZzNjD9
VefPcNVjGhp+Cw4ISrFzkc7QQv5C/w9Gzf5PoGpbO4yqd81dvbERTaAbVKs5D/X2iVeaA4LmHGVx
19QnLiCViVVM1LTFGRVyLZ/RkIv7tR6edRE9r6i3GXoY6wlxwjpm8ukTrvpOqu5iatujql4yL2Kc
S2sjmolot5cN+dGd2Q8FrMgkmQDj9S1N54GZXmHbd7L6JPMqk39VKSZv4a4raoDFjhNkf4KiQdhM
eadyG8oupmrXRVq1Qb6VnmtfnuONKOZRgz9nHh+wrnxaBq/TbnNfRGfjbavzglKbnxlnLRyX1L87
FzjwkA2OBnUCY5u3Vvy8KbKoqx0cuFobW+dhHoOQL90PLzQtr4bcVV/IkwUx31FV8AYBh3fQ+NMO
DLjygbnTlC/dhZFapHj5bKsZTGQU64Mz6RZ9HDMcRRq6+9IxayQyUSLEVUdD4TLEwzMKbfmogRY4
aS+6huDq5XaIGHY2VkIUriPrMY6StuIAbgGqWFerM04PesLQnJd10qAAaG0VF1/97VCf5jQNLPEh
4l79TspwaxonUhMRImLBpuvdoMzR9KhN6GbXNyqsk2XjYAc/flFCbn1aajmBo8z74+DsLANFdxRr
Jhq5vsKWG0MWdG54B56N8YYV6zTcOs/98ZFMl8veu8q/iWk80K/kMOGjBayoGa7viQqoZIO2UjCp
UNEoFwzYIN980NWhllci4rlpFmVPlVksMKEnoF+sMbon7LPI/IuFEsN85xCOD1D58JcX61i18u6C
AHEB8AYxLqX23rk4SNVj1qVAmt6It20+pmWZAEM6zHWPRAVKb/BrWwh9Npy1S4h7PE/MznR42/1s
v8r/XsDulkzTytNLN1f3oiCeUQQF2s66SM8IUVV63V0boA4uga7jLBACKqaaJRcA3ZXLi/4TW6Km
W6CzHtWXYwEgSuNNrB+lfw33JXvrf4k0d1Tr6XeusPDtNCb+D2+uvwadGZ4zMZYhT09N6zfoIQgs
9GphSrbkrVPdOAi8f1+MPXs0GJ9IkoVcbCLaU89aGiflOfKqSXkc8lk/mokErf4JSHCJ7UrIyKL8
W+o7BAtIIQA1iZ0Y70sGpnG0clS7Gl0AG+t5Bx4DP+jfr+yH6t52wx7mYA5t/UyTmuyrSEv8bTpt
fux6IMw9T/jO0bFsJk3/MzkVyxmHiPMWlK9o2VGPJgF/NZCpyDyvG25ZNlVaO3g+kRSzHuhc0Ap3
jDngdIMXXYuxwA7q/tvXW4NKVgzVmsap7qGZ9DXyH+zsYWQoq+ZRM37qZUgCgLFhV+ufaVK5Dt0i
OCRvz+EAf4ibUOGSQ5LLobEm4tOImexbUfTZIvcjche6aZvy7Ti0F7tZ1yQzDLx8FiE6NhXHCEp+
xMgg52e+kpL+x731MezVXOmJ0MzI0nE9yvZGJGppHxVOWZ2bcv3oV1MSSG+H7W8erhyTyQK/hy9B
ClBB0Ln2QbboR5jmsPzhvC3FcnySa7t62Oqoa2lHke5fUHFMhnkJr2U0R9w1KUHCho02nql89r1j
lURoqDyEyf8wmHWXOCqKqq8VOIOIW1g/me6/TB1uMOgG9O27PDjivvdKk+4175fKOZ0ph/JF+Q50
eUnk2+1IpMITSNvjw2dKozNPYCVPaS45lZ8WdZn1FEhczytKzXMZIm1hnl7xSDOKr4nCdmslv8Jc
MtDc1I602GeFsyDjDJ32dgqsPwnYZfja2JBBTi8gHtWh5laosd5vnBzudgDrvIDFDZLqEljWOyoI
1z/2TYUIXgi9RpyUSPYliJybysrqVQ6qFu2GSRMPF0L+FhRoE40oQ6rELx1Q7zIDjdsosPecKQOp
pDzMRM4Vuf8R8iLGmcxTU62AOdSahO4qSpFKhg9jsCRGxHTRdUbL4+QCZ3zS24XrCbcxdFmTkpvQ
Evb7guE6IXWvLRQzyLhBmqGF/4ULTYBgx35McIh41Q9zHsGBPZx5UXddVNFmATkgrnBIj4K0kY2J
H62jKqraoKOD8fmkqNZPd8k76KdV9du2oAXQYfCgHqWxZIPMHtnwnhh3bohBRVOxs1fG911RP6Ws
tTpeK45M+2yjNO4jIyMlx6HMo0B3z+yKycselXsRKpCQnVs6KMzrxuGTBuJkzr/as8qzySCraf66
gJk/sUzD5VOw8RxulxD5VIz9B4QJrIS9oa7mlS1FnheV2ftmuGjzK2cQy6QsjvnkfOGK/bHD56Ym
UOhS1bxTqti0H8iAQCOT6DgqMPA8mVUkrVcGHZamRd5Rvav7VGrI6BE22UJ33uCl/3YnDCdwyaGp
AQHG8F26M32UsQa415znrr1SAiGodE8VTWOqb8c3Yhpr+TGiJdEdVCLxXLyFuQ5hWOdMUs2HzPWK
buJoUViuqlFJbcRhiyQJEyBhkuwKkZkX32XIezvl+tvP6JFdt7sIBTyNE1JnaP6FJh2wk3B8Rxda
ZpuBDkzVc9hnX8OeoAOdFYQMMYhrey00+OZYmVe2kSGeooCIBWgH7uu7vSZm3CyLZgxkDaxHtwlW
+wkNSMCZhUKikY4NgW2C88usry7JoCuNLzx2qpE6ZlFHln1apBnwolPtaXaRFm0/9Sf1nDQfCL7t
qBm7iiUBzxPvUmYpUdRFIYU2DjHN3oFNHt+jlMId6ngcYt7rRKpaYMNaXL97mIBA8kAOc6ASQPeQ
EpYZEDQunbE9wUozsuf0KWdo5pT2NAwlQN9J93d9O75GG1bQGbfirnpNe3I6DKBEih4nM4Zv/R1C
XhephlL7G1jAkSUFtFISX/KXbUZzaNH4f2OXT5RcYrfRN88Gv9brjB06AK2vSqyeCUJR5Z4tGGwv
EprudJW+nb9jyrB+RvYRQAI9qb44iS8LfiVh3aHOLZ4IdZuWdy0z5GmOfXrdjNmbyAlkrFNnMEMv
qP9Qowms84Pk+1ZnV5o5kYa14CYIL9cZgbSRG/COo3LBA40R/hHTiJFJ6bOn+gxq6BpDbnedZnhJ
XWx9bAsTMwFqrnrryUUFYwzIw0x8z3Ak5u4BoL6yCVoRHXvHIiqbxavkiL+fxU/L0ubqbWtnS1KE
rQLrf8mUJabKenqJ+XyhgPcKxugxOAP7y0XRnnTw8DOEeJjo/DWXo2AtyQawci2sa7+IZvl9mI3/
ztmgYJf0P2lgJaIm2l2+IWxJW3kaZsTXR5B3gDeVPMjbD+5t5Ae27iDU4R0LLA2jB0uxSs4GYiSk
P7Ie224G3/KPB3knHONn43OPDQRwsO4gORyN4KP5zzESE+cxKqPHNJmpu/3mKtsS2nODNg0QR2D7
h8ep2AjECbtyJockYWYUL1gyw+59h1KFDlEo+Oo/uha5yMJGs7lPwvP9aulp149cY/EKeRfCNok4
/+OXyKOy9VbYXKQfJza24z9KhnREYbUzYeyuJWXVQWfy85lEmvrO7O7YgU0GCvf7s6Y1WM3SDEHl
Hb2JzlvCHpVNMzlS8CpYHq04yRziFDyO0+JeaNitfpFWFSrgljCMApXxY3wPzuqi+80X/wwE+5e/
lCh+ziMmCkXLGUJZM1h1vza6caIkTo+cVzdDR67f1iIbFlMMM+7p3LxC1I9gWEOlN034WmVnvSfU
gK2vK/G6xfoHV+pXYHpdVSXwFWuFsQl9dTf+WvRlrvfNjJnf55A3LjemPxXf0JgXyLlNILScrGQM
9XFzTfEDjkrmYIsVO51iCpafqZdyhXJPA/mEKJmNh0USqqNIejGozgnSuUMhGCSxFKchp7lFLTYa
CsrFGhhSPsx8MOSJFxLQp159GAoV+TeJmA7Z0CojBBwOlpZ8rek2J1ipLYzThT1eG1rL2jMsKFk8
Dp0mTL+Ctau+DfYBbyTX/IAa8tJKxSrOOIm2zUeyq8xOXEpXO+KAe4Fv1DFEj3A7EA5v61ywxo8X
5CJr/XsldJ2YnCNYWOZFtq7G0i2HuF9aajdIuGi6Fa7EHVOZo4a+TUzGUEVL7SSRRg1grNpTIoX5
Tk+YImYpA8tFAQseKNP1zwlCTYDcx5FttantoayML9yPxfNKxUkwy5UJqlnT0llGI2VVhHcd73Q9
6hBzU+8y32zjBem3TiPZjRElWHc3Yp6XBMIk3FDjGApQfa/3ohLgwRdcL7319ZfGObub5hvBq0Fh
HfoyUwq2kWFAqh3YGY8qlD3k3VdT3Sm+MUBf895SEjuwbwfPuIpH61hWg04kDXTsgCMWSFLfNzCQ
7E5sCa8MrhGhCyA4ra2RoSn2NhBGmH4QlDEBJVybR0C08uSUMUUFNVk9PPzaYb+EWxmw8C2UkA4G
HGXbav3btrf8+VP/CAYBtiNYP9Jo8RjH3ngscqy4ZhnjLL/StwYgHq6gCDSvYWxCGHc+3cviEPhJ
D+PfH4uIf0YGGa+QAOCmHH1aJYbocf15JzcEHZnmlg12T7QlLeh7ulijNkb9S8uzRYTii1K1i7KD
mfijJwu+OdNpbDOfA8ald1uagR4ssj/9ka5B/OWVTQpOeyRh743cIQA/trb2XOGoph/qzuw5mxGN
EDZrUAGp1pSxHa7zHV5BQLIiXZ+ctJ3V4fP9jgbk72wpGUWg6Qr6nzAe0WrStVLJpb2L9jUZj3T2
0LEazhUWXXAGovn9dQJmIA0JG3dBU6jz/nQTBRGlDRQ2gq18WbbGiomKC+NgIGcVrsI3Mu89tMtR
W+Eu6gxfnJs4HqCSG80GSHwSFa4M/7POWYuZvpps84GNsJf2Z/eWXPiM2rUZgso3xN9Q4fcBXUKA
Pf+w/x7KbYXl6+XUmJGpfhmiaxBXPadjCilWlz+45t0nli+sk6IjV8MdlQgMXYi3AQEYz2kq6ZiZ
WsQ9h7n23KQ0q8mMxxKR07rwsmI0nIWiCopAKRFiw12dh8qsf1uinkvMIfYiYx/eNzWIo10MrtAg
sBbMWP67E0j2JObrtvhVihrd2kUTAIMpqwrn1ieSsGJq/JsJwxSDcfw7xg6AsKXhPk369DDop3jb
dfk/PYfiuA6lUNFHJ7F1c1ZgtUYSrWS8UX6HqoyvsVoZC5T7gVO6b1/YMVgV5WSfOPNbftKcZpPf
SekYkwJnYXP7OPubk///BFIYUUURs6u7Ojv92MJ4r3Sz69iUJdqkoR9ZiqPcKEM/fo8a2LqH0GX9
scxIKZS3vbxqTeTE51/Hvk36TsArB7oNav/LRSLrOpY377rzD0qdnqvP5K6ZoM2HGUTHUX0S7qrJ
LKfQz4AhOUwsASEap5qtl8yZe/+7xTcDy19xpUVxsvrH660C70Xv6aYuHlr2hC9yQC1pedETV49L
TQNopUmX9qY6owSrpdndcxpXsNh53uLJGFolEhmCsyoNR1+RzAB8DfwuE3XTf4Nv7maRe3uo1bX7
Xpnh59HaxKYFiLmAh4s2rj/yCYrcq0W2IFEf9TU5Uyen6UgxRkr8aBYskS2U+ghkOkVdx4NqJUmq
HGMiOcv24yL5Az/uVkvdH9CGrqiP6CEWj16Wdt/WuqN9+fySUJHi5SK2YjHApy61dR9G2+jHeaIe
NZlV026fRMiWyR0lC9+mdVp08wrZD4/2iq+oBCtxrw7EiPJN8Jgy4M5Y9jioEU+uI8SAn5uMQYN5
LBW4j6p3cGedRYqcfOAXVNRxHWAzYqOKEqXot8dW4zoVx2/C3q+f4HwINB3/CQHNIh0w8/7tp6TM
TV5xSmxUweTBqIXI3SfuHluIVibipUoPh8KLYl82jnLzjMtRod8w5DqZ69L+zwIrU6vXCdNU2EBt
lIRY14Td1/ulVAYrQLyWlJC5BUlxgul9B6YZH9N2V8m3rPb1mi9ofrJB8Cuae8wThZ7wypNjv18z
WtiPx9eFOFvpIATMt4yRrIIWDp6y5TVOWwCWB3OaN5+4F86pGM6MjWe/VvbF+x2Gslh77XwdHCu9
PkuLnmJ05wHxFZgzCYRkD/OTgmG1GUb/D1Mda6243OMCdtlQg7oTr0czGRXgf8c23pZpG5e3amHX
ELMgRbpSa2RuKoysWHGYTBi9/4hw7LEcAkvx1QDYVJEPw4I08T5Q4Nu4bcSmbVt3PTxzOjPVkyqJ
dyRPl9VSdeTHGACe56IHIIQlYi6/qdg8nXOYB7D8kZ2tZN8wZeuIxLKj4zWVAxNIa1FL9dlhiLlV
61IZVa6LYaa0n2T2SczcLpZDbvPBkQ/ZmNJXhSReTqPMqX/W1YsyhqQemHUEdgpUINZGQpdOWKCT
JZ+cpkV7SWzs9mE0xS7sk9M8lGXSxMZegTstixdTFZFTS90TWEb8ejklDRD64RJbNC+gcgea/Ew7
DFX1RGv8Fr8/VrsXynyLGbIOAVxCV9zxvAr2wJMLc0ExQwtCr4IpfnFLvfpJIjLU+VKYoG4xx+vf
/9U0XinA9xzxG+QixZrXp5O/mYm8lOptHtgHtZzHcboEDnfHSBDZOgjzrt+eSFRiYWHAjda+3/sJ
Kc2H6eVTvLUjGsnzUfoGc1/KJIlfwQ/ELOwxIIkT8VJqrt9dBtRqD1vdy1ya1DNAvD3bqiHRo1Ff
XA+WfKyTvhA/rfULDNfK+FPtwk9pQe3k0QxmPOqI+YlZCs2Jo+P0SLuN1pEWeQqi3JcCZFP9HUUt
NqySzv7O+9zm8c71QyIr6hT8SmqBApWCnduiEwngwRAz8gFlfqoZ+lGtjYgI2VzXPWGlgHc9OQmY
QN4EY0hE8/dIWPaf3EynTXPK71/JI7Ep2TLcD7z9DKtUfBeb+tPxfGvcmCb6h2TxHTgGPtkJoXJM
+Lv4gUxohJSkPu+YBfwD7zFAm0NjH71KcoXHUyR3Q1Ygy/8l1tOk+8iNcYWKbBtxF7bow+zN6507
+AlI/AOAjuhfEknNxnheK5v8Rrk89PaSy/HyCrvCqzRF6RIk2p4vcsKSPZpj+yK71hz/rUPBzYim
KWtp6g7SLMlfN0cVHnu6/irP4/Dcabief4woNyfwIuu5XhrqK+cYX4MSwmCU3LIYjDiQDQ8pNCtg
TFUms9jnuuLYGq8+B5cxpxH5lnENp74vXz4BPg5Ad2af68aou10WowAiuKDTnw9pCJmwbVcd61W9
8+YEzkNQLIxYFzoQIB06F79eXG6uQQ04+arojLjnIROHiVOp8mVYhXwde+hOKs6jEWOAJEruRJn7
3IS7uqxT/BsnXkJw/WRdwMMXcfjjleZyrA+WIXxcSrde8Jy9dXSASxMaefuh3Fr/Z2+Q5NmB01ju
Raes0FBIeOG8P/1TzJDhnfdVVo/s7ofR9cdfik4uEgfKBylTylxFcjuHJmaJGnRe5CxyWJX+pPe6
LsyidrpVarCryex6rvS+YDhIw9//fBzRPLHK4dT1f2BUsAnmdj45xbVF3Y4ksxXh3Zah1zXv+srK
S5DksD3pD6yxwtJuiecoodr0JlLafrGSNDgBjfrGCmZMUA4uDv01StTo7T60zCLJalyE+pn7lT0F
TV2g8gtjckHUYXBqBknBraoZnwTqu+j+Rx3wkeAZRviBxjN30eHf9qKBwF/FlasvynVx4yMCrJQN
WktWr0u8UTyOMYswwO5nQRYRy4bJCOIMRgehS/dtBUZMm0KyET69wI1+OfE1MlZ1b+blVg5o31wv
++YHJz6JYo8oKYLkvSBfxO0PLlZPRwVYF9kMF3ZJG2XT5r20k1P0xz2WqHz1DiaDXr8NeBW8FkJl
kxvc7cr39Tf6jm85m+XgC8x1vMjeqmvP6UHPle5qufkEzMiEiNxzFuNEFZ2FdYsM7c1WdxCm3RJS
rHftomX6oz4cJ/9FZO/IkX0FWv7Kx9kr4G3mtDSkCtUVEKm8dRcX18FonRPcyN6paaMVZ0CoOr8c
BOHCja5Km2iFIeMncTYoEAJIbaFGPQZlaW/epDf6+wzAHZl5TfEGzmYD9bsyKO5U9M1YFcZDPggE
Y4c2Vh9Amln/jiCjNcFSpzEq9bvOx+jY5XckJNawC0ie3O9RGpr7Qv4jE4Cin5Vqvezm48+cE6Fj
4YxKAFI+eRu+rlsF9imufGjDl0oy3wkp6vUX4KysD8VaR3dbkp/rUM9w5h//ZB8/z3AMVbSOfzM0
oNYCvrTsk0PanDCnI9+0R3hOfB/04NIEqKNIGM17wkM4rOTbUjZnQ77FqMKNIJ3xyzMKwvsj5He+
5O18MbV3WVf4YCY0yl+WrybIEG8yvw2sKqog4MSiAzClGNZ7w8rsw92rfQz5ahiJCzcmTyD1xXGq
yDgvgZ9EopglgWfH4+U1x6VnfKhJSEDQTK0Kje5a4f/pdM1y48TOMN6qBTw+eEy6Xabjc6eWr+eT
zLq7cKOxuxvGzkTTn2/zVKZog0oZO8hscXdpcVSaJ5XuC5xgWJYZOv/KH6ZJmOYZADHCLNk/5ETK
BHFzSDMaCdR22vPsAX29HPSajbpf6WpahWhbogRTmpMgMDUCkItfExO27tYXqlQbtFuw+r1xTunb
lcmxZIsccrvxUXTlVxr/G+rFi2jgsTNwaNo3kcRskZcK0tqqDqlKvKAf90g4VW50H03KSmhdNf6S
3kNpGz4Enr/DeRLA4TH5Rb6Ecdn3NHi66eeIP20QED6Zu3AQ1x19MuwFgD4afAOcX0DB/XB5dWGD
CGjgtrXVPTEQ5Tymo1LeO0yy738Bpyn3fExd0Sq7SxX90/nLcmJ0T84JDfNR6QIgzITEvkGRu3vT
Y2JFqAsdyWcCLDW3qwN7AffZ1sJlz5319K7A88cLrFyn6UpK/tZB6csuQF64P9uILqqoi/h3Tvt/
1GapCRC11IgmVdfF+hujt5WEeNR5JdLtOrNlQKhowottgh4ZKkFwQVdJ8zbdO9RKCLKJL2KKld4d
Gigw/i8Qm8Pl2fm1GMQKIoEm6vDJim8PJ3ManNKFzySErpwTFY7WJOzXdnh5oNxeGIl7IScZArxT
G9NfYIzUK7zT0IYkv0BWDqt08Ck0DXfsm7JPb7yPYEaGLnh69nQ8LgQ0CSXgRohnuRqwxmgUASN8
zAQWVqnNv1DtnipD9L1KTLlCKHoF0VsQx7bKeJT5CnAX604Xcg/mFV8Uad9AFCg5w73z0HT3IUMw
vB27mIGZUlksCXlaLBa+z5NUU8eJpuDY3UAezFAES0f1QQ86GbXX54aLnt8INBKbey4z8mwMvBCy
a9XVf9CekEEW21kmz0lpPKrh1RAJDTD4ZPOwZnXDNeAL90Wrk8VZswnoaxY7uhCHYTssfNXD+e0h
ju1gNPUXZq4Y0mMBvTujLRjQSVnyW3BsfQzmKwpB0Q3HposXbDG9YBdPM3h6liK2kmx1GkqPG3Td
IeZwL9B6A9KUYR6A8jQGSpJyW0JLMJMPc95UghphyoKOICiBJjGvK2q6cggwszqKBY4/8x6S7T28
de/xQCTpMGK0nbgheqOjuJe9uzC0SbuU56dtCXM9lIzcHTtyAD7fej5CtNJvnAxnPGoIjP75t+yt
CBobyFdHAfkX/rYgThu89nZ0yWLOGMeATx4f8wqz4PlHQyRthB6Sv2/skbmB6C8KY0VzDzY1mXQc
z/Lyb3ifQEwhMw6nZN61CV20S6F6FVVQnJribU9t6kxn1MYVtEKVw2VUxlzRzgAH0FDFaH7ujTrQ
gbuhJ8j5NfhYPQuG2pSrOgoDDo70fb8mZpSH2vcuXezcm+rMbkQhMjpOJFGVkh5/C/UPrMAWk17W
i2NdBnFQG/j/AZC03PFxC23UhQCWo720pi03tBSk9q2W1eOKjsDVpAD9hWi7w+cMLGl4DV3RbS79
l3pQICQ8HAwBp68h3Y6dqR1ly7AYul/RqnRP9q9a0GH0XIzR2rUOY2pUIFw6Vtet2cIYnD0TnkzQ
tC01SsrrVZEArSOGSQ0rdqzPrqglZigAuB/obkfU1rLqtnxr3XsfPO3uPw8yaqmwkTxho6CWQ7yQ
qx6jnrffbUZr0CfZaHoKxFAyJFRPCN28euNO5ptCAThLAeRHnxC/EkPkaEmWCZzUlhiU2LU6+/Ce
Dwdk+4W99QSpWUh0iBR1Y8R7LYLhHLAfhfh4voqjzYfYtphoJA0czR49Hxee+jhLORgpMEn+xqEo
77esH1lyiYsxnx5TicWdRv5g0silSPNNxQOSGoPMIkLur38xRZ+aKo5TxUPDYVu4zQuEmp8kSJH/
UohXnyczeU76unPvbG63PyROqBVdTSYMYEGXeO438NG3zMlFtSFD8u9OEXlrjD3R27vVW4kKopeF
KXf0mzB58MY4wExD/AL7C3jmyOgsVRontq64oqpTn/bI3FjRtb1/9ByajOWpvuqktLqPkdOOCYAM
widdejy0lax1gb+dj11PkN4FMhVxUgSz7n/rHvkSV8aL63VWOPqvGEL0EU2zjN56ULAdIgkqUScJ
P1WEQ0g2/ELJvKehFGTgUHtPCZkl4EX+m83ZeSpVp8Ini0hJ+82RLId2zGUvl9Dhto+tw1b1Ejni
N/bik4UwREgFikyW6OguTjfoy7s3cRwpHQX/eHLfg53To5pqmc/jF2YvZsmMSFp7rnLC7tnXj3A/
x67eclF1j3/tfNVMXU1sq4ojEHWTwyj46qbwUny2DAabVlTo0iKJbeZTSr/NfOq3w4862JBonGva
43iKZROaKH0u4hPpoR50ODPZCBLVLKAdmWusFSx5GbVd5iiYmZn6czoIprgvgz8UeIGGqnBEtU5j
QT4MtijJM3ZdWTUWgcMVrDc8R41KXrEu67UoGZGz5e+APZrPuImAz57/8thNUdbZi4CL8FEevC9Y
aR2ZNVtRzUDXE6N/zT8SUPmIIe87VsKMDU8xt9RwoxcrqQLSDE5l5IfSCUn2ttTAnjmiOXQprjVX
xKLtqw3B/E1gQmbXoDMIFgmntFlx7rw2gX+XqHUqp2U3Fx7ZAcllxKtLTovxY7L3OoTYtnmd+21O
746JYkRtNbOGKDmMF28oGahb9d7+1d5Skpg0IPhLaYzOboiDnRHTXDCAFGSGKvm/lIwdvwR4t63J
gOG+18grJzd6/cKz3nCjNyQcDFel5LjI3WVg8ygBGDgAQxLA6o5+rwByngIveMixZLJh/HvQ7tXK
m84EJModuUWwwie/lsvHoGyGq+r7bMxD41SPxzi/ebKDR8ByBewtbwVkyliMwbsJGhIkh86epylg
ZboE4ugj2Tl9/RLHGD8sDBe/KwMpoeH92Q7LOmJbtkjfdBPqPuUFCdIyc4Zh2setzx9iPKBlAKWJ
2s2M+1PtubBy/tPx1HfCe8su4GYNpe0h14E1leePQlqcPTJ3dtguMch2fIVZue8cmYRdEx7tf/q9
B2yc7mnbLsHUSwXYTiHUdVX/iTJA9ABFYnFglWrrA1qoL+pJqzUYKvaD8buok5kWrTI5/CeVnFeY
PXJrcTVjPLm4VEPCPdY0cPWGFptdOwtHp+6AHcuJHceiakoypOigCA1F+UZiRsbE8iCr1fFoj3nB
Gm+f7CLTNYM2CeNSqustFSofCs2mYRdCWjVl5fjf6eGU6SEi0MY8Wn0m6jANGgL3UHMvvO+G6xc5
37Zd2/xPkbUamfNcRrjVhQhcUhaRlcyRITXTE2zZWSTesALtjz1wVWFI9lmVwUR54zwnhHyFx+3p
hZ3nnfU+t+8mS8L1IxziZTHk4dxMw99RXVmopNU/6cXPBqf7kOaEQ294eZ/bCvs00aw6kVBycvaV
32psssX8YQm4neHP8of8EFX2dnaRzgI0tg8Rqyu+j4yWl2+z8aJ7jc0HYZlnfNvP9qzOsWPmh/2t
0KYqjI5JaVj5PR1gqS9jO6uYJPMvsRNqf9iyg4CaERpQxhQGrHZVxRzsJCvuFIrSxTA3zolVB2wJ
Dm8pwtnq576J++E9f4hr8KtvFC1qJBPGDNyHmdt/tvWdx0KjI7vgeGLnjivnnzRiHhd7eSZCFGq0
5NSt12woXRPh9t2AXb6W62UC+XEGf/qkKNXwukCNvW/5U8L9/Oa2gklF5H0QipHYuf1hILP5Qk+G
6THKyx4lBR+FMEuEWBB0x86LlMT61d4XcKuRJJ1zs0RCpbQdiyW+yC5i5UOXe+DdZWWxDcohEG3d
BQzBf0KJDvdatuV/mtmtPWRJsfNmawaOVwajHj+VkcnISgbNk9BzVoUf2ryhbZ6AdCImGv1YIH6P
fu71G7c/uX1wd0WAfC9j/HDvhEPSLiV5DLZsCtpDSFV8kXMk/W/1UvXFaN3fjJi3AYJI+dpsfhNI
mhePdmMzWWv0XGAVZNpvtUuZ+GQJHgouT5EuTeNFCz5N3rBbkm1G3K9a+ouHnR2JAtQaCiN5NPmZ
dEclS9dTgfvTtVzdpwC04UCZvxj0cZnSri4dT4wiJHzfELWbe4So6ub7X/vbPcVvC6SjqbUxlAws
fA3gsSnL92JkTKO6Sw9tzbqKGzQfILwSmjo2iuSrgZfMkMakSxVHurVt+H3chtz1hSGV1PlZ+36M
pyaadczUT5tDUJzpcGDdKZNX1Zc/1Z3kGwBMDqepaRlRMGxWefP4CDa+dc5xtkcT02BfRLF/MC8C
ydegzFwNgKvBglIrY0EVgtfUzMHbjunvO/H9xZ3REeUpElz9L2U3eCRaCTnQTBHvm8jddOUzHp1Y
n8GSCoMs9cGY44lGu0lwJN4nelQhI3FlX+SXtE3sWrEk97z9Av9phrWif2fYHpKWh5F2iHlIVD8Y
kifOolJZUCN7uJ2yhiMdUWE1/wJDod7eldWGD3yfk8NituE+c0xlAQo+H7psyAUF7/kWVDbL2G8o
nf6tWsgB/tUwebzUX5U5l3Wmwwvv+es7rPCEiy5pCOokSMrafgF/5dWVg94eml5WLLptS/WWqFdj
UY+hT/4aKmaes6XxuBbK2e5aWkCtzKIONnBkyAUSkQerQc5mA3ffMjnkVNUixkqsny6kj2cOof0T
JQdHftGbxq8HMaskGB8W9VxUNcLrVPKBFqbSXV7x0vwXokgMP921/bUr8vsp7QtvnzZp5hP58Gye
UsU3pKzV1bVQOw2cbzAnSyYUAzjdFNRMjCGzyWP2iN5QqbAHOW4GbBN3w4kvKwIL6l2rQVHjPEsu
B5M8UZgeLsS69xanP9t6pUlluviqOao4o9VvMYe1ZJg5fN21K6z0ZMFLwa5Wv3eOQP+OPvJEyqC8
aCZ7Hd+XXlqGqq1+q3ppLHef1ZrlCl4c1zPC71nuuZx5Lja5M29n7kHD+daO1KNhSgIb21bv1ZRF
wxWiD4jM8cScMfsGNVmQ9GkMAP6z6KTHctiI5Ooh4yu2dGyqO+7bZZbF1Vzu8f1RqpVe2J54fvxn
nVPRG+LSSqg6j6eS6qrIjalGnlqW/XqaLfdZmpRKf/GtOFZiFMevpxMB9VRZhg1txAT+9zWYmXIA
0tzXkGJBm+y2pM1FKvHBx/oKNufleUXMAa+AqyYJmZKYclD0M7eZP1w3FQhI0hx4H0rYCfAgPRkc
gym8quHPhgMJkcX+b0huGubj2YOx9XlY7WphjalXFPd3dnXJTL2Ma8c06chwC55JFF1lGdh9vXTG
EYCbfydCwMppIIHatl+gzRl/TQBcPYF91VxwdM9aIeBPsUUpGeMfXa64RqJuxHb24A9RcBHn4cBJ
/sB+fOqkJGac7PnXQrf/S8JtH1TD3zn9c5xIRMSWh4al8YCMyjAuhJ0yhRTdg+wq7gCvvWiaH8J+
iHu4ejzKD11/bXZrgJcWiVsFkE8TOpD7y8in64FJxJhEH56BUheXrjaJDqXtzkputV8SgXusCZHA
lYIPmelriGn/uCKEagmCw2JaCIqdv/QOg9wL/Dg+1jYQFvVjJWWTK+kosV3Yh+zNqZtnINkD+y9b
9zNe4jViwKYl7GKIXNVFENzOi8/X4Lz2OGXPdT/kxb46DYCiY+bdqpwr5+015f8FvoTBNivBesYy
sN/7tnTbmWqDYwOqKb2FBpsR/tKmftzZFuj18sKBjbkKNQkos5SvNZNkPhW3ipnNgwi0h1wNACx8
9yyV13j9GWeMfY/j+v3pO66nnVi6o0sw2YTjlC7KFrBl/nOm2+eAPhm+288VzS8aOFRCC2DVMgxb
BzsUMwn3cszjiMMFffoSie+vAdmm6VrC5JU1Atg/wCDe0wIszj3OEtW2m3Atkcs8NGjFiQyFBdll
y1/FMkUUK9oB0BCusGfJtU/s1jnRDVy6f78s9k/RPXRJbFZINVx9rsmW0qYTbKJ9nMqcVh9WgjXd
7mcUK2HYCI8Qd3wH9n7nvSDR4dH5cqMxgDfhpjbxzBj6wqmxvtgqWi+yQmNEu/sBFBoJ4+U/ajBy
Hg4LAhFLhXh+rJ0ZV8OXgbLffAix7JhTfD4L6vNYGSg3Ofl4cTEm8oGYLl90l9M87+o2tpfUnppB
hSt2efNRWda3H+R82PuwNhmy1/+IdQAacUciJoT7vvnQqpepPjblwZedCpsVUXwsB1bshuys4aVy
GsQKdbggeOowCAYaDFjQDvVhlWtnK87rAgG4Qhugl/Rsb06Sxm4NrvB0VJvgEmNEAMBDc6ocxp6s
o5l8y+k1efsoR1Mp3uMRUsAP1Dla0/Rax6sCyRMErVThT3PF/azzBiPj7kQ9IN7sJUO0rl70Oje8
4XXBw/wWRu4AEfC4o6EpS/FefI+EBkV2om8YMA5dx3BLdYBgAxaml3A10QVRDr2sTnIzDn+XvFKc
SNNWcpneXJpGF1snwGp/veYMM1K6iBfwHxKHupS1TwFzSK+fJXW2iYMZNVgp+OmmRMB2MYt7N/ST
EXspj80xPvIJgvlu/y50gTloClcc/xrGCtUmBAtHIt7xE0ZXJ/fpG85u7MMuD6iDrOS8o/lYbvtI
E8/BFEiDZ/2oQDHXUI9VRuGOizwDW3Ts6j9gEhj+UQ0RG06bfjJ02BGqvcnXhDBWD9vzNemVf/Vr
W0y9jKdtsPzP6yroDnQVPGgVUngFcWNfqQQ6rskMYzh+RjdlsSIMjrE6IF9WTEM7kn2pi17cPlAo
OkcH1mucdldbxSW/x2BLr5ypTLlAdcTa323t8OrBatVO+y0azd+/TF53PL46cYLOUFSYTPwCYrrV
OzwP/HSaxGG6llkmweN8DS6A3gerWMlWprcuPwMy0b09Zx88QgrR2mAKjNSLDYEk5RD1uZKOWLFE
WGNkuvvMvaaXeUOneBANTzQj4/5WEu1RapMUqOS2driFSQn1KFWUtEWvKbGURk9Drp4TZXbMrojJ
0lJRXBLGwiV2ZV2hR/2QPr2O7HY/ehSIRmEhd6/NFLYNM7qNoIk5bq6oxAX2hETeAoJohIqHQ2pe
aKgCp/5i7P3mdL8MVs7xle86x1lWblf9HgEninueHczQRyzEaN464UkUR+E803c6bumJupiDJD/o
SnA+TlMBgq1iBi4Qh2v6z7jm3LA6X3pzgGHEOgZ3RLFyLEsR1UIVKQem+GD8VZuqepFfyCj0oHPf
c14MBjUnPQNQIXaXq6e5HhYYoFENN5YsbIBnV9JEEL11umH/f8uFARWTHQ25gATHGexyEsQWZk3H
LTRA+GMHDuMqWtm4WpEg0PU3nRcOztsnlEavcg/eT/tK1SKhWiBYD/3weY8Z/CbdCh3ha7rcK6GQ
ymWzbWnQg97by7mY+K4PBgfWNByfrBDUjYWfewVrm9AJILyPrjijgetDyUIrRQ4QQqmzGZ8GnHnF
dyKy6WKIQnIHSOhbsbdbAX7xY7lOo6z/JJsvN3kJC5dwWBKiYvIu8dJucpOy+tJFU9YWb3GIeE0j
cE/mpYZsJcdbiR/YdGIFEdrwLW5cx3auW+Cbw8+Z6FX+BikPWphuHG6CewMnncXkpNGpZoiNK7r8
52j4/PneiagQ7XmalYNDkR6qWP2eZ09Sscl9db4WMd4ysX7G946Ft0Q3hsZntvB/NDxTLhZh9/pj
Tr2MBDrNP2X6a7KTsPBEpLdtYHmieOdQLnth22etkvktawpN/DFamG6oe4wbDwWWwbuqilaxCq5H
SUx9ccgKSyZz9oiWIwbNHHlIfvmE8JprQJB58tswIUl15N2X4wZiW4EV6p7zOUBdSQMTeimJpplA
f9HCOXhTI4ghY4LZP25k+yspkgLnR+xftd39FGlCAkx4v2hK6hvAlAuzrDq2HJHryNopIhYzWMgT
sJr/jf7HIBqE6cgsJ7ejo6CJsCdeWhQowC1tseE90ZITdIz9CMFiKzsy6yiCerfRPz0zwGNmQ12+
/bOgjtEyqIPNzzxCcm2FDA//cN2MjFj+DgMVc/1w7ckMCAihoX3NtRj/oSUW4sIFXPl/WrrkOjBH
1BX5MsmrmAmWmNC7kdpeTodAOG9BogtWde8khMTgKFY3VODHG/6uj1sB2ngZabSxNibAZ/ouJA6r
rZ7qMEEdnDB9nMXIo22nABsPRsF3oLyP0xTw8mjMtnsdPm0D1h8OashECS2xhPcMzciQizbGl2Bm
e3Eyh0YVQrCk+3OjRyQRFk4LyLHK+teFIBpCifb0YEe7GKHWUxhuwfup3kjs3uh9Si2pu2gTo7T2
AZCmxqgVwqzZrmWhEptxPLYSVSCSwT4fIAOr2tHZmJkxVAgRMWGVuSYLweCbXcEq+x+9hYG0jo6k
3Vn7RAR2O17qdElZwe3F6nwDzH7UlVW1RuiUV8FSbYKD7qckNmgAGbCP7phxGmnQdcvCwhJc+Ppb
lhQi5JRrx++nGWSjLB8ToFzE7Iryg0hB5iTAsxA9SlBacmaRjAySOX5qQL3Mr/koRaLKW1fQwded
H3UmwL5jMPH2JPdXsrFUDn3OiQmMD0AJdeqCmqTNC/Ez8dtWmce+w83zpg2Vb73DWeXLEHVBMRpK
Q70PM7l3oVukAIDLuvdOk4mjie4XOutyTI7oUlVqLXfzI86xl8seWj9pcMPWQf35c9ahc89k6YtV
3/qzasFRKGr4XwOjDFq58DmeEx61WJM4Uy9yligOVvOJOuS+UR1SA/f9NI65B7bVEmEbA8kaHkw2
cqWkF8ODIgVrtDRo2stz4jG2x33NHkG9QUjasww3q7kIjyltvOgKHgl5xJ9m/n9Fk7rvUCdlHVdN
4jEoFRoTzST8K4tck6WDJoVJlwXr3E3EfcVO0snB+EIADzvhSqYLeSaJVhLwMe6F/DBcFVth3/uO
Bx8PCGEpPpdWFb7vGk5gmxI8YEqeWzswzZwti70J6gdr1WToPFP/vYylhiUEfgB1GZuqswcyypUS
u7+3LsWGnOHDGbrqO8Pg0WudIFfql+t+3GsGVu3mb88G24JuLq7QSKefGMB9nXww5t646W4AmJ4h
gyPEk/DGADWo4JPzP7h7ZgmfvyAb5l527+lYOetcKaEvTrHSns/sIvQyo+wK3iCA9mu+ksifYDZp
dYN7s/R3mzlshTNvpuJcilxtZ0oh137Vz1W8b53WlixnPdBY2PK+iJEmME+1/9KC67wwFDdCqiZm
LzPwfZmcU9sSG8Cli1Kj+gze0Q56AmBhJl6Jz4xuYqchb7F1cQkMLkfu9L4tKpT6wBB6jKwZFq69
XgYD1y7FM+InXXAPD8WwaJx8YyeWBJg9bME/erFGQl3sV/y1TeSTlTxrWAdO/US44w9emdlFvvp2
HfQk21dL+Yj+j0Y5yyqClqIrxwX9KQa/xeEOnAVsBkoM2M6LocBK5QNu8g3dQg9L7LOjaXy4XJK9
Fw7rifxG9sq2WULrGLOGH1jOZ2NB2E4AWyziKl9ba4IWSTLu8EoZah1nZOlMQur5d5sTii9c+bYA
hRy1Hxe9yOhiswjSR4zqumkduVT/NI5jNkPMpJfnYzrErCp6EAhSLBaXyp6i9RZ4oRHtov5ax+GD
KvOpMvKN4cbXWoAUMPvZawoUt9yp9ybnzzV1XJBXvqK2b5RH5OEDg/a/fMuWWaQbEW8I4lzsLOWC
NXrhKMMuBjmyn0fn9UrCXgSbHy+Oo6udUbpxHLuKA6MxIXnMEqkUAIC5CZNW1STgJiickLnwafLk
JyqSy4WQkcynLbx8mLN21lWR+aQ98wJQRnUwqJ/aRchO2ERzmc+CxPNc7rINRzsSvF6nVkSF0/df
hUuYaCoNDnvih70sIyhyYtQDZibHnVZiTRfovTYQmsfDGxZ1QUVzLBqolLybLng7igXMLLi5zwZT
oQY7ui5vooeuWg1jV7l4sKmCKZyimqoynwnbW1NG7Laf5pySOzyeReWCT32FbMdIFbQgct04A1/g
Qo2ic1DUyCBUVR4eIMS4fPMWAgaoCxXnLZ7jQWb9aCnw8sleV9riOMeYu4UXpKCQ9Px4DLzyw4M+
0t1XXa7C5YvX/GMpSSRnAZzgj2TEq7S5AZp98re4nZ5Ud+oqERZuZD1+/9LN8vmxE+6VqVUj7gL8
F1acIpOaFJowHU0qyXBqqa7bQAtQoe5lPW9Ax8IpVRcJ8Fy+YyS9MPk1hV+o8mbneoXd6FLtvhMl
Ql5pE5cZB8WBg2K+nyV1EH89p8WvN4w9D3sXhY+tJHAusjiWqXIxd4lIcdGfA8AHmCeJ99j9EvTl
PPYPI00AFCRkje2vEt6S+9kAVGceEF7JDmu06Avez44YwBjdoIARQTkz2LbMR6gCcH/wtSHaUUz5
hY5GPk+oepoElFxWAFINWmXFKHcKOxAhcd50MuGb+tVBVVBXGleOgeLzBRhuCgcEHOrOVkc8F3Oa
cDxCEsYx8lvSSvzELcjj3n0J6kSIcXMeFs/Ft/XlNNlsS551sqsVGXxFlzPwV9JazrhOfv5T958k
DcFwcEDsdU7VrsZ/8dDPRw9z9CHhGwSuvj+rymPHPRuRwVJdeeYBwdB5QvNoA49684Ic2/75lU7t
FrcXvf54ecP5UcQgoeQHe8nX046BTgtVr5FLS3mmBGuQY4zYKVLVjfyuCwQ9mlH4dS6KGpUojIxn
YHcAop1/sl7nE2U53JQ2NVxxI1PSgDpS0G0gRMcoWevcLVLQ2m/lx3ppqpiB3tkaealcVopUhLfd
di/FH2GkyCOyNomRX5dbJqqsJKduIHAAhAmBuM4LrF7kkCzenmjaN9gAGD3zIKXXerlr1smZPbCX
BfVEXzXd/+ZbGG6RjuAFpUqxYMaiC4GWEBzB7ApuLwXU2NHP0xpBJe8KR1CXq+mh+mmN5cB9afgb
fGkDmfC1J0xGCSGez6GwhWWxZDz7nef5F92GGxzij/Gqxx9VPT5amLdPZOS1WzIsfTh1cYmiA8rM
XgMWMWzt/cFlI+COqYKTcXnH/BMCnd6sSRZnJThSoXC8W943n27jsCqNLYg9D3HS/4oEWUwMEkTq
nLifVBiUttgGqw8uplEsAUErcsT/kM7n55Cp49H6i8euuEdKti7qLiVqHfVBn6VNqEysLMQRQw78
PdLslPzZkTbfJ/fplZ9CZWC/ASut8hiSHeX2ANNGYZgeG+86kOknS/DGR0HbFEm8YC5NjkYzOpaS
o7wVTG+IsqUB0jbzQbrNNg8AMg9R9omlPe3VX3B7UC9SI9IRdBQfhneOdygcX4rTR5B+u7p24g86
XfjCziOmEosGf7L+amAZe48RKF2Nw015uA/gXcOHHoMV8BGPn02fdUP+uRqNlogKsJzzHvp+I0WN
8lFdQNDs83mOb7FOSFxvKAA1N2AIRzvrg7+rK/tEtdwVSdq8wrstwcr0bpPvlcP9rVlcqKuv5eYx
HQW4K1wj9pk1nS5//rLyPtpppOSo4lzFyA7faEIJ+SoFeUKSe9RACzE/iNof+GY12BVQXkpbRWW7
8HOJKK4sTDchf4WDuAIlxA0JjS0ZhG/97o+aGkD5SUYwge80zv+A0Qpxa4KtTnLVoqqxt1HGrBwf
8CKA+Nb41fxveif8q3DY9VGMa4WOprngzjecEwmZcCzHwp2/lurQSyGxvXmRpN7z/a6ehv+zFy5Z
cCm2oujPmJJThacfRFvcBsp7jvOSzk+JPI+amRCqIh91CZ2OY30o9NqoyJ5V2fL9L4vH8l7StXkp
3RgzIa732KK/j0ZPazRpXKAISSdFnrKhI8SU1JDLJ2ZoPgMgm8pArTjkLa7348i5nnClv+d/vdfN
uSro/rES9Pts0wcIsg+lqFP4TwqDlsb7xC7oHfncBFYCfeWx3+vWYJlBDqjQ8rxVqKsHYnp/+NCA
rv5A0Eu9Ktk3kXCqlllDZsYS82eENXg65rkZI3N+rBPMBWAVbhS0ivuELycVg0afHwmcokKnbuA/
56RoYCug7sh97XOEnfmJo/KZV735wKkn/9yNdaNTh4n7MSoqwWPg/S46HilZBqfuEgOoPzL8ppp+
YMejs65rTDaQY9YCfPZcDlJ7fByyvV0qEpuuRnZv8QhJitU0Wyjn7zQP4LuJNY9BE1TYGqDazS1Z
bnr8EnnEB/nEpnRa7BaXMd4BKvvmAxOqCSr8cfSz/V6U/wcCDgC8h8WcJaMLXffEwDf4Ft9WiCRJ
JBxJ6CwTLWyJiC+oo+h4zCldTqtnJjk6Sb/Mnlj/d+dSH++SAmGKTZgtWy2o7vBBY6Cs+jGqf+Q5
QQoVlScIpP+VPSqMGSw8dcfsAvP8jh1BYfNal8MHHBnQx5jMehtUIGux8vjdZpcwPngSGpn7g5Zn
VAaScBcYOimKVEhJfwq4VR6tBEchpq6PPUbdlS8s84iOklaabrhx14yhJ7i5Sapj1y8jGzFiSU4q
+f7iRR5qymYgcBv+hgEHWgTKsMEp499hdKYLmWziOcIk9N1WzNZoOteGfOXJxlcsz35HZoXI8Q98
RmPXuSg+pyZhCrMBZo2eeemJd76NEvCjFBDWq7Xm077zSrrX3OpIqkAYsnr+7UvPh93RPoyeoUgL
jGJVoKO8dtvjGjwjTMKULlHBAHG5FxXphd+8lHjHz02Btf+maM2/mPDTO2meb0zX0wnVoA88ClVq
x5haoDX592+t6UOSk5GfV8/PIWgZNpL3LrA4cfvBYaHucN5Fy+29QI+R7zw2CkSDrFfw7B/CyCe4
hgwKVT++FxaBS1tDm95vODuaJL7plkH/CBOraW8ArwZr9BFyi/yVrsn2aZVL6ddZoUF46yWhSsfy
fPQygoWJDVHrD7FQkEg6dHb0r2ZFsIzPq4p3Uj2yIq6UuX5Cu8nzNb7O9v/Yfidxbvm2n9MDkm1o
hsVJf0URUyG9awkbPSEE5UieMt9XRaTdVP2GwmBxqAk06sfjgho0c6JbNjj8Ee4ZBWqwZ0ZPUZ1y
Ibl0Ms2HouVkFohbDvDEvWxB4xRIZJWJPnSMtFyAsXRLajx76rOwFqiWdqDFtcD05nmtX8ALzHuX
Rpnjfz80eevugCt11b0V9V3Gw24jZ9kOKF8WjHKoZQ5ko/M6uNvdgH/62uTXNPm3+p6WkuPuT8sI
RdGQrzx88Q/2ow1ffJgf9WwlkQfCCDoxmrQ2Y6r64pfGrgYPaBY2HRXam+VyJZ7cprwyKFtZiFDF
ZmTDc5VcCixSeSTJDhLjeYDKWeyQR3W1IC+20qX6FhifI8YvFKRHhrCyulH95g+EUtk0TIyOoWQl
e/po8eRZ1eLbUggmqq9/occJEzpLNeMGLHgXSEWz64ym8roliT3TiGcqudCKD+/0UxX9DrDPngQc
ZGRRdSytijUAd1YrXWQp0R9Xg5MGFVPZR3Sc1FFe7gIPOMSZvmOg0GMu3aX7I7+gm01p4qxgnq18
NmD2oiGDZuLsyE1dAH4aYh3NxvZUhd8y0kMiPV69Qb0Fz4sf+vcdLxgdGwS1XteB0nlWOnFBvfZO
3VCfdo35G++99z85rfrXnf30T7+is3R6q/7lX9fHuqeEm5nF6YPrl85Y6HYaEflxDxracQUhiqfW
I578RK/zKSwEk77yJY0JilO0FvAaGIcxsj5D7d8bOdlQ5UWni+qxUiJCqqJ1Um2EjOIIpgsrRY8+
MT0t2RQwQhaDsqsVSdrge6Cq6wtear9g/QEcjB73jbSslRk/5XXiCbPU31yRZnZZkkjPHwKr5wPO
xotjNu51VZFyaZ5JCVtOCYKLH2AT5uSeLQKK/7Kb93qyAX2QMVHX5q+jxGVlC/J4PCqrlHKezBue
jnvg62dCeoHqTIqymz9X+uaNw9TA02NupimXVY5Bw6Ofho0OVwZQ9ItERDmJhQoFXLcj6PiquOJX
8tdPZfQVJU5EhuM+FXIeKG9Q/OyvX7J6vEV2xmHS9LWjKT0BsJoJv51+BxD9Rd+22TEN+XVGF9eL
x2D3pIl2/+692IHJBiPI1QYM65ENSuL4gL5OkdItj9GL9dI5Ryb+ieC1QxF9o93VA9S8cGczJ5v1
7owkJtZhFC/T0yK2cNGO1BrY3QuzQAIu+rTupy32pS4YcTBtw9NPLpg11aoBbDiOk0kFVgSMMPRL
r0rKWUQk3YDU/pRRtzy4+jALlgONFwQrTpHY7KAczsV3rHefx24rgD0x5P7pO/uzvoou9YmvtGk8
lk2TWQJQq1fARtB044bE/HkqE/qIhVIBxxDnVBpGW9Vj4CJArnToTwg2Q76F5Wpf3r6MXw8KbltK
5X098vZ2oVVRI1m+ZmDSqQsHJowYKNtKG6Qft8ClYPAIt8NNLULMYx2yEve9PdpAFkv+cKv85kd4
R6A78lRayDDwqDLJFyWJ+ZgSvEBOXR4d6nLs300KFXcFYPhENygEEYE2Um2TF+q4V/i4m8MITsil
cVNh6og1UBI3DlMxJBfiPcyeiIgxuirTovUsQwZz+SpcShXh66JCl/qLkTX1Ghe1M+L45W1CPXAt
tBG8pIQ5BUfKCCrrEHxYRqZnCNy+U60AMwxcjdB+fuObz2pb7hWtUZwV5+s47HFYLjl3m3yXXFV9
Mp0S2XSBSH4Bi+Mc+ZuouQzgqBCAp8MEn6x8EueIx1d2gCX8z+bK1vRTVgjroLE5HLXoLo3UsnzB
xPYNrnqEj5r3Y6u2zBzsMRs07hJQNS7qxeIjo44T1el9g7sbYjDq3BLzKYSVa/JvfUhYnVR2ZdVG
4S+b9i1M/o0l9LBRYroe3GrGF+d/z/pq07LblYRRStKsbmVr2Ul0gvPZZBnI4FP4wcg5e1LWXXbo
o/FaAVTclIEDGyKzmlRe1GBDGxqWmOjan8+2LzbeR+mVZcobqbt/jhKNrXmAtG1uqcWJdPMqI5ym
KY4J7naDt7tr2lmJrO5c1lrz+k1LvFwAMBdt6H4XIJCYdu0dY634AMYm7wlIHrghNDOEZz59ez6P
Qo6AjYPm/ET5j6qHuO1pJOfXFSvQkOeBrtQ3ub1e7saL0EsvbbBg/tTRDydjV6xd8c6KKxnfIblb
wud/lkelv+4OHrs3tqu+ksUlSLK8aEsQCB+2q5E6LYSvXy+u3LpaubMFzm751EmooZCBCAfHP73K
JzD0Z8OcIuwbvZI9SOARrDEAjqGrCvIpLJQXPAxKeXcLG6x0qM37+zO2b/SASK7x3rqISpWIz05u
3H8wM4Dt6CcNB7ddsTp0fSJTcgv/RaXoen9hBP+XiwjdNBxT0f1bU2+xffCg+boW9AtklJKPa032
QQ8M+dJd12RURVtD2ScBhD5ryM+RU2oMZFF0Naixv/p4BgGT9t3pX8f+LT3LUXKsHlAqt66+nRH0
GhchvcbFETCleKQaPmO6NlnS7nNHSh82L4ocegf4IHXMxHFl67no59BlwAUKCWu8JJIRWiWfcwic
s0Lx1jiksum6eZL8bLAWZZ9P8ugb0pzi5KfO42hrLJZVUeJNPEposE3jgrZ1oDReSfGL/LO1n8ti
n39MrTMVlrYvBUruVCdFjEGjALXs1BqqrY7TH9dZG2SLQ0s7H8dTjtQUKIgF2r6JqKbky3iK1qiE
Atw6s7GyVZne2t+CiC84huhP/A+hQO1DBtBS6LFk5sRdkcGRkS3L6owDZBxda8iggcaR1IXfk1sp
WAa8Z6/TtC+1qb2Xd+dJhTYhBp8biak/x+Jwqivv+onA0fEGLBuplZiCoX+7s1pYRj2Cb/Je2O9c
jtaQbSoyKrWpHC34UyimAxjIGUTQeEmlC799ZQ0NTv8MVdIfPinKBBOH+sFKEDKJF1qKvPeVFnoC
ox0EjfOgk2ZLZzD1HysmHGpfzNTKSunchaLS04SXMjMoZD23r/Q6QzVzRSxeywweIutgHptd0u0M
epovmOxqksIqR1vThXdqPVzsXFubZ9tKOOol732eJMUulgepo4t0A5lyRmwgSQl2dtOwDf/0IStj
cSV6sRl60Ldhs44a570YpWagDrMk+K0gCfJlCYKqB6DjYRfshu4z8sOy4w4GXVZALXeFDrgzCAKl
7HIENkTutwNskOhL7qRFIR8HKtm6PBTRd5vI2sS3Z1ImayH5i4jd/qAFHwLYz/PaW3Fv3JQy40mw
WsUdYPOVlmeaDxKlBdky/BGZTCOke4qogS+SAMHAgcDoY7hcu4xz4B453ow1GD8d446fmv1x+3mV
lzGi1gqGeG6tVdzi1HRsqDV7ovb/1wSoexXOnH9ExTHpOXEFwRofANgBa2ytwy58ytQalIVZbmc1
dt0cfKt7aMn0h1YNtDbntyVlqqP//l98hOYSEe1ouCnN6SD21ke53MBBhlOndKTTl+MF1wvmYeNK
9Df92i82kw9hLJh9VgAaHShljqtIC7Dc9GYiRPwL/j2BEKeSI5bH2lwJV0ytJ+y+VIEzRKN8peWd
fmfUKIZH7Dt0E642qnSIh7oHW7/l+/5R1zD/bHXz4SJg7gyy3Mau/V8l1oethvTFw5REbJ/CC9MV
p5ssyqxJPr8S9btzTCk7PhGT7x9sRJa5Ill0hiGEq7QHSIvJciTP3vUBiE+7gGEFDghWi/XJqaaY
H3XYG3Vu1ipKO7lwXy6xUCsExHDU4cZJ5zIXSmRcGROaUdn01j+MWFabXyHgvcdM7zwvYItQMa4h
gBQ8D1T5TPLNaC3z9ohTHXFV20A1BkkVga6FOzVoG+JRCEvVvtpRK1KN11Phk9AIdhntl5qDooBG
ZPhCNOhtBqsKWh1bBVgoB9bYRdHJHGQYKSqbxMtyxxoMHlbFNPx0vLr5lsCGdPZmgfu4tH0NcYxz
L9jz6oa796/Ur24Dy0xMkCYxfhcF0MZ7Vnejl+t/CGkANxtBJ9qtLqgIyyy+Dos0ZSwINBxquyEo
u4A5MdCAYnHHvAEtkll80EvkFOseHebYKvRvROLvQ3ALeLLVa6cOCx9QgMqbBh8fchhEmyDE6Ixj
KJ5QWOY8RA80pdCJSpMuURvD8ZyfmkeBtefn8KfhM2pVYHz8oMabJDhXhRFF5wUpBi/giwEtE7bE
mO4QBewsSHfRWUpIjm8S3QU6GvLWZmtUwEF+DS7XX/nmXkSeiQLmqGHU9Ij9YFJOaKnTY992QHzB
QsCJ425h1Nmk5siK6kGJn/iAn7hbRIIwKOgSCX8htz5/pgKqp1/RPKfys77oIbHgo2SY+gW+gbtj
ZS3B8JHKv74lI2nbquRmlyFBT0mh12O/O02RPuWJRC8rqtzxUyzpVVSbEyLKyQY6GSGCg3j1bpzR
R4aP5l3LQo3YGw5rp8ETZuSp6A09MRDl2ZUExKPhurrjTDPzGAAIhgO3wCV7V/KXCiY9Lcd76fZ1
8XnPWgVJKcB4p0idh+nWKKtmKMDEN3098USsAJGuEd3uW/J6fQx2DpXhgQB7i94/8HWKXwXMVpNi
xAVTvVApu9/Tz6xBsWU+xWOxioV7t4hvl9ehEH47cEfnkFt5OQXxQ5JDUg0442ESXfOsKwKENgq2
shh2q3GDCVkrL8oL65RgMHdWTaNct1slJyel7cfBuE9uGBKqtqYonyjSIviVpvqQ8CbV3ZCkdmiP
+45PAOlZzMT8hNYuRQ8OCMJ8PZf2m8zJIHejycBK8K4uT3U7TbdgCTORsTjqgRiwPueA+0tNnizY
RI0JS4xqkkxgOYsPG44HixhwwDr/OR9b+65cfcRERhSC0PBRq7lpdEmOwbyBeheUEzDF0Pf/nTmT
Gn6k3tK/No4OdX7a4tEHMr8Gh5wmiERru9B0C/UhbauS8+GF91XkXBykjHfS+MY93xhAOskU5DRG
z+JmXQnAJKHvU1l039uZXH41zH+dxH+YuubzGyv6hncsQDOqYS7iyo9YTHz5H1ueQ5xVcntRWgXv
kDEjTVrPvvt9MIcvx5/ke16rPCm+o3J+hE6Zi/rn/pTDFGqm603JolcbEhzFxFD/MS/NBwDNSIbc
09Gd4jeghZfbvfRq9XAyb0bMWbD1d8OsrFF7LREnHMCwcePm6khRXBrWhwZP31/EkwZVEg8DNP34
LGKI14WD29kxfOLcpOYvK6hb2Aga1NT7onkbUchdO4JalOULSgKgCVmw8BoAZ81+C6wZBwwqVCKq
4rKfB5Gzccu04GtLakaT7g0gy6MpGrYBpL5JPWozCwZEs2re2Pp1wgkaOFAD2znyJZCErCDJzJqU
PASZWzebksHMsbB5PubgwmUZxXcICHJwwso99mJFj7OBMwK/42lgTCePOM9sZMjbBOM3UqboH2Xn
MSpxLuDJq8TX0ItyGtxdAZeSnL7pemsqvHXgwBIUSp2YpF/6FGz2oHKKIXmm9kNleAl9wk66MPzY
evq3orVQieiU+2ioeCHI6qxVbgYOke8dnQXVHDb5+D5VLd14bo+eX50Fuj5T6q+QsyHmV+ghYekM
kdXuBYM+Z0zj9n7PDTbjJFphmUuoJRdjBJ9g1I46TSTBb70Dus6hMxEM+iLOSXCq4sc4KjJUDaz1
3fxDAGgfgCH8cbErex5EGq8sts96hJgztKsAlO8fjCbjhz45ch2SKnFy1dqqp6fBaN/lWBO9I6JY
N9GBPnnNN8fr4eZGK9qTuNLZVMlZNIoJt9kAAw6ba+onM09/lCjaKBm2jtbdhHQT4/7HdmB1W5BH
g3IvSOipR8IaF3YIVncUvAfhTzKCKg1j95fm85vxaEZvdR2bzna/E5IiPNxL9Fih9it2YZ6zS2Dy
A+PuPQKjDDypJaXKNnYD2RjVHOUFARkPhpZYHsmBhdgsDD4aWZOLrTI4Yt5CbaXUSQPg15vuxMFt
I9RUOZ0ZPPDEs2FhZmlmGJm0YxfR9Xs7dZJpJ7+orF2XSSis47XzL4wH2NyQ2i0EyOZRTRMbvGIz
Oxf6YHF0R0rymT7FhJeLdxb5ipqslUV0VWjGb6SOHMfSxBWQ7alNtxrlR3cPRzEQKfj10+OgMGkB
W49Pg8dBF8E/Uu0E+QUoVtvLwy7EXxGIYC863WIGRg0cBTXSTZg1AEeNnl9bfy3sAi4hmdUBUzaY
kxUyt9qJsO6QJkIBF+Kz7EhQdwRDLV+z0SHfE9SAVHWqm3C8EPCYn8AUU8PuFrbX9h5BIc1VQ3NF
gYvZ4ebNVQQGQIjm/ENZGyKmRecezxiAbrSWnY9Br6VVkHK4i0z501gv4FSGaAT5GGbq7sWqAbj4
oY9mH15hdNnVSonW7m8a51/AzfmhcaZP1v6MDIOZ/O13OG2mAuRoDzINaqhCCuiVeOEUtRY9B23U
EN49FJdTp5+MI8oONbYIO5D1PosSrkBRwHU4hM8HcT8bO/bNN9a5TIWhe4uQmyNYigvniG7LGNCq
anJ6p1gzleONrE+NEpH8iamTW4qhc8S4gkrTNbas7CI5uypZx1bMJ+2NCowq10roalL6RB63hhTq
djk/NEkEb8n0tmfaj5/PPwruK3STcs1F5XurUlIEryiSk+OaoqAty7mJKvngy9pFU6nlIl5dUsas
28PKuwgSyOW44x6qDB3aFq87AnMe/81ja9SgFs0+gFSexk7262xyaonEPc49EfBPJbvLQIVmKxgJ
dA4etsiycP+qq2ITnby/P5wghN44I3VNAHcUNlSyyLkUKvILbJ/OqubHwF+bKyr3HVJL+ZNOCxbe
TqvgffnpRTl1AhlMLiNYLDcjwJ/GY2hzSdgMbFCUUIUIta+5dbnn8RueA21kdXEJNSBVdpuNv8GL
tvSLWV0aVH+o5C+D8InMf/KsA9FBHFS6GoBIlL8Jv9RjzzB7G6s6RBBBP2qGe9ps/Rs7PDF4G5rK
TLrkFuWr5ZiEe4qH+HwXdB/Ixn5UJXDhhbOg8HWRQDKYNmV2u7h1+TrOnxZXiVu0PzsP4runNgxJ
wNb4s3Xq4cyOKRY2UvR2+8pg3UkMyc5FO2qbyrsxuLODZkUDlN8ZPJ3HMdXz4fbgARaDoNyfnmgK
52RHsEvs9pbR8Eu5rdCDvmBTFprQCU/z6Un72J9D5IBjGH8BQ5fJnfnk+iIJSyxX43V5UmqTAVf6
QGvDqDbdqx5K+DfRAv7PdBXF5HvMpY+EX5t426nsYQ6/3tstPDOcL9jFGj3Da2Gf+J1aC4XNv0LC
kfy/Njet2cMs4hBznFTchNqgQsUNG9fbQEKjmzqQ8kEAhxma9xvH7AR4YW7Ifxr1T37+Y58drojM
nSDer5tK/SWtVBxLzVcutMMVafVhY+cy+zcW+7w8CBjEDHAeWqquPcFCf7Fd/rBvUuIz2jH8SBvm
wghnWLhPo8jJmgjRyMeM3CLmU4O296md7bit+b73rx5k60NMlplCnFpQgiXhafl+SD3M/cO4tZqK
+I21lDuQW3zhCbsuZ3fi4aQhvXroRSckPERDiqR4JM66vzK8HR6/Zt2B/Zn/7dXAhYM4HHj1lrcs
uj5wF98S6UcA8gGTIO9GPiM7jnfj7IAhVC4IjcPmvi3J+YbIMxCwMFgzCxJTTq3Sq+eaCJ081Iie
nrtXZ70XPk8Kj6sMCyhPzLX+dzfdOzoYu5MViFVu7yEAQPJehLncUYVdjqqoYeaz3VkTwtqKTDiC
PQJ1PhPhAWYaZKjh7zpb49Ih7bTgnA3P3YaK7Zxgr1bsTWZSjGZ3rAXM+J83Ovw6oRvQN8o48Pic
AgoGlxptN2EYS+eHIa0UJi10woUbP7Wz8GHvmy9DUtICmoMsQNLYgBSxXgewU4FrYQ5w2Gc/9brN
rNP/jy4/oBo+jbCCo6smyQln9rLME2AXmUu8Te1gyrFsQr26wxJRYFSZmyMiUsyhNR+GFCKQVrBa
xfPM8VVdAflRmoZ8Iw2qrQOtxl/d5wVwsY5tUvCd7yvvmiP5sp6c/KL09cbljCXJZVeIha/6ovwX
resXXnxvzKi3McOTkBXGQjY+jSIzGnh3boWKodz3dHaeQzx28BCi+kXOKInDMW9AvmaxVtJQCkir
FdDBRFBMsF92T7hZs5iDfM6EAIb7MN5a3FKkgY9JRpXvvqxBd2Kj0hOmDTTVtOaVZ2g8EIt5E+Ht
ui8L0EP3d38QKWBst8lzsy1HKoN8E3gk89dabxBiHLPgg4FTxPslDL+/Y6wt9BShDVmZrJznnYpZ
qjol9MMJ+gV7+GeEP7ef++loBmVpF7nLKK+4IXcmk2PVwImWd7koh8EQ1wCLTkYJaZXhuuBWZR+/
6+TkVVv76GAhF27MsnpoNVA/EOFZOufj9CeXaODhRSo32i3l91GQWBkULe+i67FTvSjx9gPOnZcx
paHWwZYMqsWFzkCax+RBWhJ4+F/yADuDEfj6hZuoQVai0vG6uMRusqF7ETdfykLjemeEqN87zbxZ
SQ6WA4fLjoIVvEI9yWd6dG6VXoy9EJTyKqK8+Nd7/jf4AYR3WoKmE4TUl6qu9h8WGaypj6rMkNeB
Qts92J111JDeDsq8iis6wNzN/qqnDuufxhgp6sw+YwncYRIbtI8ZJFSjteQ7g7UYpnepUrz2Rtkh
TaL2l5BG/t70VoTcsd6nT6ECRNF+xPn+KEB4CJbjb+EDn48H9UcC7CtPXxIn7yp/cHSwGfVCHAAD
Ug3GkQuhkArsqCfumnKt8JOtM4Fe2ne+AUkw7d9oryZdKSCkqhshqP49ORM2E9zlcMMB3h95yc9Z
etf7HcA6y5e8jCc3NZ48M3QQsF2YdCzfNfiCXSjW1EQ9fdU4NAVvh1MiTuDBRlki04EeOfx2IYB8
O9AWtP50clMjuD2LxLeKzktc8LxgIq60x1OoQGKwLhqFUxLN3uFatJODRYFGYDtZOArdMfSl85Nx
iATi4WYk/zhXDEFM6p0DyirfP+OHiyT6UJCZUzEZIyWN69YUlPJrGx1sWaC9r1ycQBrjCRw15RCn
FPlRLa2UhqntzCcL7563UNuneU5tjn1Ehk++wrHnHMcTzYQm59j55OwLIfSn5/Rp5QxDrlhY5w2r
Drlh4PLbkW6tbLnHMJ0ajApGBbjxnNqZ6iyNC46l3OAly+FWs8DndmwKNXWH5jIoROGAqKC1ak6K
gTn/YWl9bGdkdl/lRLpJmTyslin2FQsPF3CwlVnbovl+2ws6fUtUKBAwbTNiqz+P9a0MAOEgPGPd
6hTgO89gCYNhbYgBTMBZViUv6AEEaq4G8+jsy4hLRkGNlEsfpceYHKNXYJk5y2+RzXOl+jKlcSbK
ItH5980J6W/nfqrzGb+UY9R2jLcac0CNwbw+jeAaEUkty3I0Fx2wqsbsWy8uEhhh8LJoY5b3heKe
bnMVtzfa4Sni0ZuxR3XzP+/576PGpHN51HQBX04+IiDKh+waBh78P2PnZ6PTYwlFaJvyoLt+Tpi5
DxiEpwKgLnhYL1zEZ9z+DmjNWM55oepOryXtjL3bHb7ktqK4gO5JGk8rNUSQJOwikHZToek8n8lE
RSIMEn07Edaik9TI7NpnOKdjXpYELX+XLLD2gOU6khR6wD4FwR2ImIf258qMqt/bQJVg3TlDGB/H
uZ+6xkbjri3NMA3oh0bZlAog7KcZHGyjcR0njhNhlNfGE2v4xRv+xbDRVAq+q4wTOgzEhauV021V
GPXdiYQU5TGltlR0bKZylxPiMD1VQOTLdj+6ir1sqMFu/XAocoiK4hi/lWK9i4sbOyj9dpBx1QX3
byJq+VHxsmvT0LG8qX5WqD03bhbW0m1bbe7B1TrvI7JWIHGTwh0DIokFBxI3j0bFttLNFexI26hk
XuQSkOZzuIlg63DsUhjsyiffOmjnrSqo8igwtdM49gg/xVhNcvl6vauv+4wZGnceeVlR2EWLHkmg
BP93wurQ7vlFiMAFpeC2slDjHbnJsPdvAIy3fcqOSyq+yh2+XdWigv+bk0xD9+J5fvYYJhk9QMwJ
2TA78pP9pyHiqvWK6xkBXY33cpqUG/0FNERzQC6bm33Qu4wXgt3Nw1VNQ9jDFLrM7zNO61Jw11Ef
bGVL+01yjTA31r5yRUbsuVHnj1rrJ4yYzPuUEhCTzixXyP7g+VxO6aSuFyIy8w27DeV9D//hWtYO
BB+0ws5QZdXTmIX0YOOvTWkvUJV1FSRRl07LB0FrdADfOpJPwRFSCKrXX0qf5a6EqRw1wohpyKp8
SBcw/55B4fHofC3oqxZXEjkQ/ykZGtX9RY3LvsFZe7F3TAANhLD7vAs4Ns0CtsdQQw/hfMXc76T7
jVrKjXT5MBaZfQjurYMeiwkJ8WQgVbVmmL3BRdgANi85Z+LCi6+B3ZgT2nVhqZak8IWo2D63WSU2
A4zvJew0KrlmpUjQwJls2+pyXtLzH0SOUGYY/IwUno0ypYnEPqtanSSi7Z8TLf0zAewn3gtxHQ3Z
NBBM08ePw6hwwmbmbCWMgUY0/+v85jorAAIzaOOtgwd/q9JSgtf1/0g42nJRNU4esP+Ce+S2muk9
sD4J4RehU9P1Zm56iFwEwetl+ghbMlwTO3e+flVx16zYVapj4ViAvfvwN12DpunS5vccokS6wFzI
S++73dn1ENXzc+L5R9T7bEcRNFLVdFA2Z+yjzrGdMP5SIyRhsv/69XbZX76jPIrF0pBJrjeCJUEC
poGGrr9TNngpZOOZBWcHp7ui/nlfgSZsnpXW5LYzOr25y25YlUxOBBxQk0nblYf7aDWQIC1FFMYP
sNbcG5vRNJLwY9ORqzhD8tGBtWDfqfuILPSUTa+R3qiD0HX73Hapa4kxaOKo4UzaK36NHxybI0tY
3fqz28rLCO+TDNEpgn2QAUep9bU8I5dBLuZhpwSr+rlnKPUZr2VbnnWnKB/8+bCNgEyKTHLtk4JF
l/pJUQca4Kr7t4KV1mwuyZLD0YjzuIhP0ADrtf7dvDsoh3mlw8Z2+MNMD9oV8SdUAO8HoO3wmOV8
nF0C/zdJXc+4CGlg9X7eopVC2srDY/gcnVbWt32nGoKPzVgJkbzgvpM2UG7gm3/sLQZZsGiP/lCB
mIP2ATmsdPVntpdBiMo0peaZn7RoFJoZf4MlSW/8abq48iyZvsaj18P2ebchRDP47lPIB+ZZRauw
+3RqUFJ5T4jDijA0R8BswjM2ehktS71tLZDKnCoIvIzYlwsRPHDQzvXCdwO9Ox1XaVU3EpT7J71l
n5BgJtOrsfYvFjIhf3w0X0VsDb5oI+Xp1acIX9tJdh8UwEkfdan74OFmHbFCOfi0tM+NcyjNtDQT
UCnFA7Ci8D2qDKz0Y1oXYO8VzCeFVdqDlZbcbFkwwHrrw4NHsk3PC4Ow5WwtY6Y9j1uZWqmOT0Tr
slhHy7c3nhf9MMexa1QBu9vHmZG+sNMIEIJ5cwhe9/dvoqoGuh7U7Mh1KkevCxAtGV8yA6Q5WQJ+
iapRPg+9uM+8HObYKkX2UPmEeVWvo+ZVBnxRUiUOOrfrojabhUpT7eR/QoBpgvxyhZ6ukQAvUlxE
kkA8TEXPn6WH79zcMew8v/cy9hdWxRL4JZ7i7Qf+K4m63SHa3jSbrXVUnlMjduAW8beSnClrtSkh
mZC3DtGRIZDxqITXEjpVNci4RboGW+BYAweD+uxTUocGWfUJv34Z/AQob38PjVUbBLwX9YO2dHCc
9BR3fA+piirvoVgM7GgQFIf3ImJi/QF0aCuHRbWYo9GOudKiauSwfTa2NiM3WEW9qnWO1uKIvfqF
a7qQtmKz2F/GHvKAtrVrDoEcBjV9Bilo+n7qGyOLNtMOxulIY4CcuvvhFCpS8vKq7ep5+DJfkz8g
sw9/kzaUqnc27Lv9/UMM0bY0BVmnXmC95BasRpQ9Pvus/X+abBx+Q8N04YkYh7uap9yZaJrj0UWj
ZFvu0NOxGTm4G9Jb+QESa+2Q1QyJTS2rM/3W8AcJeQT3TiSRBH9lEf4RyUk6UDlkTuLv46/9sL3s
hToXUo8isHnYImD6fqrWajaijD0wbzdSj8tcp/Ttiv5KpqA/cEt1IyaW+8hdo2F90OhxBUUR/1tq
A/6cj6FZY4hXHl4HLQZIGAGKZEER4LmmvCjCnK7o9qwoKOAo5f2I9a58jMyneaPMFD4GSV4ffnmU
ItiTRW5Csh914kdLN3j3NtA46iVGXBgtAsvB+6sCvcv9u1FdpkhXHm/Mhzp4LkLCsZIOdeX2ASoB
lyZ2fwdfPk4e0c+8XVKkYSMC0VUTm9+MCTPwF95TWwMZK/+xSQHkYMU14asPDQwQYD/Kj1yY7YBk
Wkfkm2AFgEfPyiPQdvl1Rf4OL9WXLgeeawChG5wUPUvJhW41SQmxOz3KzCsfnzuO/bjsOlJ80XwR
lwVOPFKCrINUysvk6gzavUEdBjXI4mpl0RFIi6mPbGd/A2RCGc98medv58JABKngGtvc0KrNrSGQ
nRN5Ua/69Lcr6w/xd7DvduDQvm5fTD/Y2RzIv0FOL0uI4HDpnPvC0m4bE67VIalTEWHsP7CDPZHP
khtIvDRpjF1mBEJ6ILINjqj+EUghqwj3DNJuoTUxrNgFBM2RS/pMciRRycOq1QxM8W25iJqSAhEn
QOKO/ZkeLV2RHVaTt4SWHjU50hIM1kbiFGGaU7tXDDdNTSFkVxeYwRYagfihlpojComzlDRWPS5C
V3nOfbckY/ViBj03NqjpYUZNPnUpsduOVj8hM9w+6duW05GFVvNG++Qx99mc9KsEFpE45+fgMfjm
6gMGWpPqzNjxvy82oCRTXUlnCwhrYWA+j5LdwFf7GJAul5s9GOyHgDskNXI15FZ16PS1VL0JpIo2
lmapclnYBbJ+cJ5wd4L/LJYp6NE4oT6Ll1UvTptQOv33oJVya9zu7uFu8FB9GZ8Zq2e3geT6AnHf
LUnGeOH6K9CjQawn11jpl3cow3BWD+C+BZbxK6dTKAELSvY3+6LYRM90AN4Yji7C90EEVwJkanta
9eLDK/DrpfXcUWaQ6yHALF0GtN7P/Ku9FCRhC6YgtFL7MJjF9x3xgXUj19pwBJFxr1IL1G+Gq/As
YKMkeA6/0vWuz80W0nvbIJvhA6TLZxLdUPK92hNXQdoJzU5dmCv5XNJbU0qOCvBukjtGtesrdUXQ
2VwiSsflP/dqkv/rkPPRduQdCuLcfBJVR04Hrc1VepUuKLpOinS6p5zHc1plja0CLhYasFhmxrCp
VvbXekD3iDL5pdvM3yn6tS8CKp3ovnhElUdH6LPco3b6NKIpTgMgjX4a4MA2HGVFTYNTNYyk9hTn
4kuNvaId9Ei9j5gapkU6aUZ181n5beFMu8xcRvCWw8WokoHmK69Bz+YcWOKAiFeHCSN9czKrJzxY
B6j2A/d5Lq5x/EFHimVOb7MG0B5rnUH9G5PoYA08I6GA/r/BkHevGM5g58rJRJCY1VjBIQQvL9WO
JozmLwjgRzrh04VovUX9Fq7GXn3zBia5uLDbe0aoDfLQS/mnQjAJIbrQovMcaj647xy1ub7IQS1C
D5M/IwbEtj4FQHAQZ7sVbRtt7ohXRBVcp1jArJ2batzJCJSlUVmxqMy3s+v+AgX9WJqpzIjtFf24
X0Ok9S30pWyqLDIXh26r14GyA84chabmieK0HwaJ3dL9leL8QTspzjkWBpQ5xZy4AlC5+g8XLUMJ
H95wqhx6MqzNezkTfUEXHn/TXc6vEdD7FZKG6BGSS0J6mGH2aMimrJsB2CPgxg06l2XLaXc7CdYV
FKFp1e5KN6fZImYVvK4oG1i5nErWhZaxtxbgpX72XVi2glzLHbWMJGvw/hlQCueInMhPUuSjhFxE
F2d2p/80vD5jHn+NX0GF1f2unZAN2WVjstPwplBKIkLyjDgD3Bn9eWhE8RVMCSw4ME26e84VMHD1
P1bM7wJu/glpVgzAqD1AiVd0wdY8WNOsEkL5ahNoyqXuEaZyYXFiUpV7raUQv5iU7YazhKIgKxe6
yq3ZgrzB9ztYrZzcbM+MM7Dht00tUdimgspAzFVpkGo33KvytFLphsYk/GPZFFg5Bdtzq10QdlTG
NlkxN7wKiwAd7OtAo50yKKLqF/L4+MtGbq9vLl4VWcOVTRgAdiAJ3+ljL/o2fm3ifNXKC4ZQtUSi
XVpZH//OnggHxGkHCulZpwxSBMI2lqFc9FW45fsdcN/40gW9Gz2QzwIDLGMg0srgnjfH5xePMbAi
vSwX4AufeEKEHM9gHdk+1lQCX80TrxgjEit960qktMoEbwLV2nROyCj+IymRyu3vsq7JcLiXbubP
BsptWa+JJ00Ir1B7LfpPvwC8giS2z7ohWlvp5m6nH4e4L+VOjlHSPalrRfw/vDst5IDiscD7kG9Y
IPBOegJMyFv5AmQow6TflujEfCpeaNFKwDzW5gwbCuuYc6WUbf5tpmeUFP4LmdMTYK9P4Scyd1SG
5sCcOJWJn6Q72HwPMhezCLSLsNDFCsPYptXfqqsidH75UxBxqldy4WJFHepmCU+C95XIzzNIi9xs
hNahpK2qyDvuvGyI1+I7aEUHHHfQ2wfEIAIGQQOmzgTXrH6aJAI7n9/ZevZCDtBse+0mnKcnbXhH
VmfakIxE7wqNGEBl3GKH9DsLmlG+2cQ+WUuxnsEXlOidcMeXdexqfRBM8pxlrN5Iv3ZMPNyBKRMR
ydWjcGsLuEnK168MTQxrAxVYulN0Wk41nU2l5j9k9i637Mh+Y4oahPPwzNvUklBLwmyXVVZ60PKL
4kpWOxFBnOsHIBW2cmhtfH3VnSSiMVh4QLvjaQzpzCEq8tqfdbgbqXCdVtPpyB/oQMfoD+z0eX1l
Jrx2WRbiok20twwMOfNu7Wqo1rNGDAh24OPcrA29xaglMyegbPzPhm4S7mBA8tj3IynPrRaZlgCF
LYtCMGNxdHMOHDQIqq1yqLU95ZHD7EAiLjgDJ0LeSuqJOKBGUpGmbzdQLhradtL1kSZOb/9tK70g
K/jGAFl3eikFzryYCifIHQwh5CgubvuJPkaHYfjb429n+YsP54v2dcdiebCgDJYkaOgOPKZqSuZU
Je3YH76vHpFP0nMB0fnt4+3pyP5qVQAeApYZgJv3UA2yXJvd75JZ8j1EM/Hv/S2bFA0OudP0Mnmg
hHIzhJ82Whwb+iJwrevnECKM6bAb5o141cvNjOnJkTVNC9stwxd1XobB9zlNhTPoQ55csLeSfOs/
dDqfk3h0j0Ymlss+XrLRuBiaDUwHEOK5D+PXBp76gIrPclENOSosQlNWDNGHxv2VqKDJruq0i5Nt
74Zb+3uPjgo8iGugAk64Dof6JcK2YWSuL2Mt8iCfqZkw7YpA8ylyQ8YQ2TdMAwUlUKg/cJ5lKJdS
zNbbgHmsJUT9l2puy2PGKuOhsVqbSkHJ5zX/Oi1SB40roB+hxcPu7We8DOiXzGtsMMtYcxy+vpwk
Mvt7fuwxViMOIvlFvhtJjO9pq8ohbhzmMVJaq9Jr09jQaXVSat0LynI5fj9SusHPQ5XHiQA+G0UE
cZDy/CZTyNIAKdscw+mG+ud4se1JcT1yyKdyPmnWgfomDH6nQt1d9HcPnjfDfDRrS10YdNOWW+x1
ZynBSiB21h8/aV+ercM1o56+Zgz4DfyM6IVNYitechJGbyr182xtl5Dh7WUf0Njf07pTPQMTCEJX
k/+PpJS6jQguxB0jnXBifOLgnULbFmXx2f+OfOaxgEbjX5ArKpycGtygnDDXku2k4BXLYtdAaJrK
CBQR2WUYXNMPjvj4Ts9R3wLvHuUufzVmYJ/ASvAsYnCKX9RSncfW81QbfO6ouIwqIqOnIslNp0QY
iNtFxAYh6ami8XCHE3JElEJzp7LtN/GWAfunBD/h2Iogzz2MZd+cJzGBS2EAtnxLQC+lsOTjW9ix
prTkKOxL8pBGtKLcI/FXkmD/LU++j2JJydZqb5d9PHMvXbRTbkIKY5NPcWWBxCiClIBgNGqdqoH4
Blx5H1SKuQqpHruvTpl9dmh0RXLtjNSyqvmLZmbI5o0RSgtdJUNtZMU0n9W1OWg242w5xWGabuih
GA5zmLCOizyN5rLLGykYM5YOZ4gDNGVUS77fZtFR54mFdnm1vd6S0Xt6zuQmXm+pVr7Ke+hxsFLY
anC0zweHKxvfe0EXqQ2wtvU4unxJGlv3bky5HPC2iZ9inTKubQWJQmF/aZRKNdfxnB6qjgnpgJGf
CS8F+pPW6TyZJ+4eJ/8NVjdMgpZtIz5ENBEHfC+nb4qcU3uljhKOktAHjWMEVVeYxzsQy+pnHryg
IwEMqnNKcgLveC7GZMe0VTyEUssWcc2O+9DmF9rakAXjEi7wis0nUIWSolPu27Az/hDedC6NG5D6
SHPR89dwHEMYGbpK4s+TZNHC/e4hQHE273Pjr2eHpYlxHQ6sBq4rityOY+SF04ma2diYaz9apMgR
UvsV/RTlaHMakI11sDdRGY8O641VINXer7lYqjKCpEKXidCEB2eW9wxj/18Z+N6iJDKtuO8WE7nG
t+IEfVnmfi/RbXekNZ9RsFJjBemyfZXexAuVEaU5r4jV9wZPuXrj4a++CPgpx/kmFSPYidAGZl7m
gyYNlxs2FVz1eoIc/dMlpbrmwoLaJXW4oZDwCOstp1ptrJClWG6Al5N501wjHrirFa3TzSGQYg4A
WGlWJ/d/nhRcdByQ7AalrNhOv9EfHZf2GvqBg5BNbJkseQZgIKgUDT6yBtbW6J4ukdhckgbYlDyh
YJknl7ImZ7fdz6Hj8dBHkUARaxsqcUEUqiWKdSLejtexwEbY8Zz7Ir7I5vQmieU7Qw73vv0K0p9b
Dk5c+NzALVoiOh/BS36SHJyrypeSclNoT9YpVP+Kt/tKdpyFdXzwAyruJNZNoeZHNzTtBLcyBEDM
TdngEGzT1Ktg7/vjWfUzUR/NzrF5XnvTLG2De9RNhZwc50Ad1ENDHLu3J/LyDviUkoBT9/1UijFN
+dsFqqz+2k/rpYngAPgdzbK0SBcS009c/U50izG9OS+ZNjbXby/F0JkrQrU0v23Ern+e1aAWb7np
VY2X6J22aFIX2TzpQv0PIXc5tI+fJ+ZAj+5tlH2I+k1y635+z9UN83Y1sC5PoVx5wGWEBzsZCij+
tNRCumwm73eUyPkCl/gy+JjH31okALYUOAMs87bZSBlqsC2xc890A3xl33taOhzJnhkJl+hQZjC5
wRT2a54/F7ukbRvn+FilVXsRT7C2/9lI5lvkLqclvYwkte+zaQ3GXpCxtBJMmM+vb0+mYWs2WFnn
QzFu7oSrKIdKyrk229Pil7QMOn7pYfTeiPi1QrCbgN8/Xmsa2d/4xyHVbtHmNzjdtXu6jHj2540F
22NzHbVjnX6xROBxMVzL9/VKp45u8qCKYBVQkatmXTQsbHMArNAMj2tt2ESi21itg2Qbt/wax2i4
MjCxQfq5qPuwiIP5sGXqJJT3v7SkYCT8OKhhRafGohlpM8oCctuvdfFxObIxjLdl8wUKYzvg9ggY
2F71R0SMoCA42jW2aO+GjKW3agPEBhnIsLFvFKYDeVm9/VeKyPYTs79OJed+5QT9T6Z65ZJ+x/8Z
ujoTw0qMJqZgaZjEGPoaXEEU5t9ax8lsRIy0JTOcGQP/8jC0xme2cmeCXpenu5i+xlCgW3e6EJs9
OimWh9PIs8agc9J9puWNlXjMMhtI5Tm5HjHWDp6dp5W3fY36GX+aRi+lk1UFGIBcXds+q35WOXdw
t72OvC4pQwUbXwCbrmu0syLxIZdzT/QNg99GqZGo85b0kKs8/w/xzxWMud3TKJ05cl4UfoP56dyI
oN+ed7qPuolfowOR9Gfo/3TFm6dH1CPee4ZtBSyY1acNw2J5bJVqDWkBTepICUXjlfuUO/e+7ewD
awhmke4HwA7yuSeFlveG44bIjPLJk2jPBQAHxkViQHFEEbMtyd8MHNOqov4Z+nCVf8odAoCemgwI
uWQ4buYr6m0IaBx10etj9gtjdeCIxMDJmeC3/oqr/NWrCNiWOHLMAQxTY79PHccx66RdnzZzqEcM
0xVKA5BzGDdQfQB5vpqX2FMQs5NlWDCqNPwLDKA6T2AQ6UbjzRtLZOCZVmKmUEXMHqj7HYpVTnXG
gvZmiPASSTGWUkVz1ewH1Ceya+p/py+cSq0Gc9yFZwewqKJH3iWiGc++FyrOS9nM2fMz+Yn5Ibub
3UfLlRA4j4TFpjOYt9kC40NoyD+gsn60DVdUfrPbjCaAfPmS+8CmbcAO5V1r8w+PGiTjg/VGCFb2
HB1/i3UboNyWee7LeXG0HZ8W1RroGZFb/JtytwKc4Qy7inLt1KqGzrHeHNiD+S5eOzKHzBxQUC/x
nJGu9ydKIVSLMW8yAwpYzoC68/noor1l3aaJ9/wTjFXloFK+RE6QHwMXJIHMAsNx0UwOD/je8KWt
q7XLdxSIgZBxF/a4Al05qf4HIqv1c3ngUdwp1sUOK4WgI3/t9PUyMtblwm2WXmEFF6sFd5/VC13x
YNX2e1f3tufqIWhuSfgMFiouYR1uLb/oSE7wQaQwjVr4KYJhnI/C4sl7Ql7uNJ4taGzzwUKLRnCO
EzIa/5W19SoFSiqneNj5sQWIUabfyj80g35qLhtE4E3F1B7xBiyD55/33v9KlXXzf6Gj41RpMhqW
joP4wcVgeQDtwvOYBpqIjaqIzYdblSq9MvsPJC4UsMfvd0M0+R6AUB2DpZgSQRgDRUhRTKZS0nrF
ta7W3GKwGdvzjQkFrbRCXtq1EnsZQx6lL0BAdF9eU+YqEHpdf3YtjCS5x1g+N5AvAWsVrGyat5HY
ItFKMbdkKJL6yp0BdpNpS7i0oXgXXbxM7aXltxzlLg5YUOKEoli6RqSCt4VmWoCpB4rp7oxK/j6h
LHR7B9yxPTCERiuBLWdDdDv8QDVat6S6qLigfXcRV+geESSATdpOiOMp9bL02FZDZUAO2tqedjnh
qd69+p9ojsH5ZGxPSu/jzkqFVGG2LcCXBNg+IN5cJRomjnIx3xpeLqUOqVVorbiZh3/cfVWDYNGY
lJuKt55wpThFdNNMGldF6w97VV620cPgY35VHVn52CES/WTYJq8F9ei3HczIpjeIuLwKjO8NqfHw
GiPINd4d3HsaMqaaAP/76CrlJW7ibA3o+kgwfGUhkRXXbaG3ZTPS60HIECYXE1BOJvVo+cFTy3bj
bFgOH3vnD9jQhqPgbDGywDHfu17HuvxHIim9zpA/Hggjxy5FaB893SB2tvIv33IUrzCpmG/77FJB
yKjSWWklmTkjwq4Bm4QHpBS3AAanl6HQmjbLeMMxjdT+iwEpNk/4uDCPsCAJa5YuhCKa9Q/mju+Q
i10OectQY+lGJFU9+pBDbP7/9QJzee63GnTXkbhqkeisEedTCitLG92xcg3YHoOeETBDFq8YUUcv
iL9RgMgvl7l9LViUdWD40pkIzabQW8QiOQLb8G16f/d1B4KhRFXEEA/dxyaQEIwPrfPW62F06Tdp
v7gp0pQgBOZEgisg4miV+Lx0Rv3Y24n/YTdxw2dv18sXCLePkmuIDd/diR4DWsmo34fA4dDV4lC/
MRx/YJx/WJ1ZSn31CrV6U/YoSXB/ZlYSlT+bgaQ1eTjGN5W4e8imZAfYlLjHMlAE9q5ZcfRk1d3z
lD80yGVuJQ3dMV+z5jmNkZNms37Vs7NaLK/dJ15GpqE251cEju8NO00Au8G/l3IaKN67nljCr4/L
wxSbqOZ7InPnL+RbJKhpCYt+X3C7DVQAJK9E/XomxrhYL2iZ7fve9T/oSdU/ctUbrZqjqdjW1sUu
0uiAu+ORINrMc02LT0TUHG+Tb0d9v6/yXN9WqERcFd0uLKrcOXLfPrg3omoWD3D3OpbtL3cnigZI
uCpDTsxQa53S4SbAfitgrHAE04+qGu/gIboLyYMCULF2C7Wb3M/uTRcAQQIVO3Hw5FQVuv2pCX5Q
Gn1KXvRu093/1StztodsZgLkaqSTV1wznFCGWGrgT+AVESyAGjRdhXjp1ZL7sKc/AiZclThKWnE4
Pa8uFVW20xmKXSezOyKs4Fs4XooQ48jGYFuKGEvMviUvRxzw3M4fhJEKS0hiWHFts+ypYRUHMVsI
J4LGauKvccQlyV4tU1G/kjgWJlwllTkZ1sD2dMX4tbsWl+Y4gzoCLgsklwR/MvPbZhftOYt7VOiZ
jXfZwyntdsAWr/EXbB66ecOuRMYE7uGPIvdQiXbgV59U9AXfAqYyIjPAUMfcHnJO9kIQQ1O4DL4X
+WszBJJC+qq7SMQcHNpQJWmDeVt0Li78raiClqTHTe/xkCTIhCbZb2g/Wi9/UAvP9V9TJ6c6YkNc
oftnNKygbu5oTRsuNSlTV8WSES908ox7kWh/hlCTjFBNv8cyPDbTGC8vGk3BWQOrL6/Fv6Q0HHoe
37oqlDbHkAPSILOKcRwsc/kcApJ2Fzl2o9Z8tVQWLbAbEnvP71+4EPdL3JulGSKABBApSrKBr9Iv
9n+1H4D9k9kRInRoSA0ANjOmimr3WJu6klTTc3ye2CU6+unvfpU32djIcs8TIHd7h0cWxwrGNVue
1xWI+W/8SaeiNrwPaTXOpUA365G2c3igSb3buE0EjyJH2qjGCi3KDPn4tAz8d3402nup3Cuvlp9z
HkXqF1Jkio0unk390Mr84ti3Y6X0A0n3SSpri0BApflxmr3+ZLUD+3CNtuZYbvj0AEAI+10rDq2U
lmXT/idLh+RNRttG89g8LNExavlVG94ju2c3A/9F4grSivtPiiS29egYsh+1sDeMtvd8aypQ9nQf
QvUYjnUI4LwblX2v8P72vD04N55cRu+n0uXKy3fNXk9M7UjSdk7zM6sU1vEgWpqh5rEJUqhgzRwK
lPCZc9Dr8I+oMyxUXaKAzGGhaPUFusy9wrroZ+uiXvS960J1GyfDb3EXe0YzcRUFgaSz7yKxDX+Z
f0j1ZQJS7JSIF6awopOjy9ZKQU2R6WQrZH8U6/koOisIkcs5M/ZRG5cg+Um5HA5ENrkr8UcrQRPd
f6xQcqDTN57Q/0GhaCjqy9hmAzt9djGj8MJQpda9B3YWsl0/Bz0Ffd7JyoiiS8OKX6xCtuPsHRuR
94Saz/RMZCZvM9z9MlM9om5TqS68ZLEsKhzTRNZnoexkaiinu/EymqXFILL30QfFhoos/bZoMVyb
9vTqDXOgYDUoVq6H/MmJrYtcqHzz4RSzFXsFOI+9/3hJBmIqypvJYCMWOoEEpsm3E2nZA8L0eBoA
/3tp0kQdN4mx0KpJwnG9k/DVvdvfNbyJ0NtAhOM6RkBAjolLiimgW9K64gZhqzm8/ihf5RgxubgH
djgs9ptkrUVk3KKZpgPXVkpNwc2DHysyz5AxyJa8ZPAai6s4KAsROHEri8kSBGFxLgMoRbNZWj0i
W/H93XAGgZOmYN6OX6Jy0Y/dvXt4i642tb/H2pEY98DPso1xONaHzTw0EHCjzvVHpuHTHzwAFjzT
pgx0upX+DPY0DqVcl+rZ6YMvplBrPclSfxP5lYDTcECFiTKhhgUucTS3cEd1MPZBNeLGn3DL7GpW
YvHzA003ZVRI6dEOJVmAcIQSfB8qXUwT03XbQ7FGp14DO7MMZvrLj+TgSjcAVcAa0dAlQ6SsAvdf
G9BRERt03utn0AIVfPZYaX8ymTBEEAGTXuQojE4T/dxHxw8rsoXGYv1BDTWvOvogNhlrlGWExpPx
/ME21y2NvFhlYoyThn6ju9FPjBaD4XSMkULWAU6rUy0sbTiQ7/b/auEhNIlK4JyO+Sp79oNRTavI
oVzZyBwWz8I+4aeMqc985hPyDw/lvln5EzRcm4WkxqRyOAm99q/r9wPqgbK5GgVLGQYKZtzMRnV7
W1dUp4/nFYk0IDTL4Y53eOsbzG/Mv1AfEOB1AihG2zSt3C95bTqC+1cRti0deAqj4tcNvXZekugN
I/kN53u6jb0A9b9HlPllheG7QSm5CdYRt/pSd/7NSBaxDj3EQYez4rShLWeNs35AmIzMaroZp+Zz
AOwm5oOjl7poCryunSop1Sm7lMhnUssY4MUHQ6tWXk0Edv18lzeR2+u0pMq3V1aCYhU0V2cRfWnv
G1hAH3dEv01C9kz8htJ/mYj5R82a9nUDbwbTP23J+IcmVhzflOjbTn+iW8WOUAfpUBSzud4xWfOl
EoStaXg2lpp1wD7SV2xesnDzTTjQJVuPBbn000vooftBnoDiN41Mn09J9f9fy3Aqgefy0r6QIkgk
iLM4a5JppidtB9cKA1OxISrS3FCF3u2+PVTrEQaUF3en7LizTZdZLCIGIDn3o99EcAjUKv1T7Ji3
KEMxJmw7TvtFZHSxVd4Tu43y/VDSRH4dyhc7X4hvv3iAncvCeZdHCmv5J/hleDpzniATuTIAjqrq
raCaQMyzxlY0e+3YUnJnO74iNvQLMpvqp+by2pC6gf2J0I9Q3EGO4vD4FJFWDKX7wOo6Bf5MkTvT
gqIqjq1CoFOYVp9LI5HEyK5xlg9CQ04TKAxQrj9d7QU8GXAfUlewKq1WfY8k3h2j+l72VNxOIfDj
AuZpQb/8vnDH4Mi+UV0Wu2Z0WctPDDsY9Dv1KfmTLN8jAjup6MaTaZsVZsM8lujB4uJRrRWj854R
QVVcf3i4638wFDs567dKGsdbfef2gPn1giSsLU6aoAWxtcNWMrNO0fD28mzXfGmmOyQIxdVSNgpX
dR4Xmex67Z5sjNheVmFDy1UcNyRkIxrwITenaXeBhGav3Sxv7/WqdWBCwe3e/qjsq1nnm9hpNRB7
e78dISIiEeqjojdbpeIptM98BuH+LjJUmnqvJxtQ1lzXb4Un9R9tSBkOG26+r07cg3tp3NYpEl5O
K7V8KSNHRJoge1bVeX0Rp3vQ+p9jZqi1Bqr+vx+YkJwbhWi3YxXoyMSUtND0tCBTXQjsv0/tzznG
bw1THT0eC49DcCI99x9XE9QTQmilgsQ1uH+pHGMDarl//5S+kW1HKpx2exgieNNyRY1+RFq1I6MS
FHmK0hrcWZWT8v7dDVkMxMpZs7QfJ/9Udoz41LMelVMYDMxuedMMdiUAAC3xjjhIy+j98Sjnd0QT
JYwHFn2h9dOEmcavfFvqD2ot/36d3zhye6IXI81npp/hWVmtm8WqGppEPL3QZ4rWPInfjiFDGDy9
OumqSBAyMKHA2dTSQaj/NrGkWIUhOC12rARsAZIIEES6PzyvylP+4BC7q9gIMBv7Os4I9lb7dFOt
szgMzPkMuLoxjJE/P1+pkGvjF3hDQfwU5gnqqSB/jk8CVRvTm6VVW+MJKt0+5drqYCc+Bc2PyWTq
w3x1kPkg+okcrWGB7UwC+DeiTro3Jo2pOyK4QFcjnJxRQd/3LkWRO76gVFrsVqXNuLScxNgOegVQ
L744YGiYJvxYF9Vp4M43dH/Wa2AIl/Cyv+mNwchquLdJCbBPW8XRBhTFN1r2kKerDrxX/doFZOnz
ExXH56Wb6ZN2/LM5s5VCFyuYBqtgFsDPrbSwZCWiPW9cwPVeJAhNHHmCmYabzyxfe4FWfj6T081d
R66/h2e1IUo5SEyzQSuskkIWT0OizHHB7CMUeioLUuKQIs/2d92i/uleW+NEIhwNEaZ5Vy4vLh1b
MHegEHLG4FJcHLUJQibFSmJM55xeTdJ1nYcD3YaIaROpLMLzTuho9Kx4njXVcRdUTbyd2S+3acGT
QmQT/tCkHRdySIaU54Lver9NKgiqeNdgAtMjVp10l05INbisUgaaj76xGRhr23lFE/xdx55LHWhQ
BQNGmrKx9OSeSIij5DHYTYBvU3/kreu3dGsrD5yWWyt4SZQtcP2fWdgpJVLChJUviA2yJ2G7bCPs
alymXUVjL8/j37pH2e3oOCjI5sdaXHymA8rPFRLwXEMmTikXYjYdTyxnicc/c3xcxn5rq4AOwbV+
xJ5vZgseDDiS/T20l1kjVi5BA6H0DvcazM2xSOoHNSeGweU7Q+mX1j6ydVk2qMAnlGqPtfzuwb7K
83ZpJyWuO/zgEFW1kEHG+e0fWBVf0XzUwDv4W7w2BMW0HlcSQaTNgweZ5BvlQr9pWjNUPdkw7qgi
r6eom46HWo3nHaUmaRX1f+HciMhP2MK/+4deCdjNfgsYYnJfjjcj0flI0pzSR+NZLTht9us+1ska
DzMa7JMNoJ7IB3gQNZqJ+oJNCeHA6g7LsIGkEAV8Sm8dghrr3pJUfTmTkunwwsIrZzwpj1d8wE56
LdDpWNfqpPb6vDDW3w0w8D95OX3Jqncq0qaoww/JENhWIXZc92fqKuc4BKUq0XJojM0csZ7mudyg
k8J5D1WuNyvi7Q5ZY7dhBaZXtVkkNzQ+SntUguv4ZEt4hXAt5+sPRcsZ3jYesnKjssqOt+fIGTzT
6kVgGzakvyGCRR6jd9FRTpc+OG5YGy2tTBOBNpKfNOntbiHe7dG1qcEMFAZHL4TJ6NUI4YXX5bNg
quQYN/py1yzdAqxpbCKPQfQtmTVw2g8wgV70RHQtJ9Da5n1hbFgIBr/aetF+3zDk0PNjVHB6d5FZ
14STTIybE+qmsbn23q3yN21Du0fBhVy+XEaAN8U4JKh2t3FzQaN6GKgsjMTjAaJrRL2RBXRDBuY7
XiQxtIqhkJxPai7S+C5gaw8SEdL2of3RhNz9+rqkMohQ7ASl3s1/a/5sPDvamIUUkJD0XsELiIbQ
EBOsTZJ7zs8S/x4Vffo7PyCVWwXy3GvsFvP87W8u4nrkV0B/3U4t8W4pY+rcgnIuqNMbns72MMh5
ltxvWWhYXLHJYAtr4nw8iCXnnFZVpYWGtY99/IAuMxBxo5ukRtGeRvLAZ289ZGdOvtPtpwcltF2b
uFglA3CmaG+lCz0DuDiamkdK67fayey+KkMIzxR+fs0jKqUPpBOdbAhMVNFBRGLWeb4Ih50nHp9U
78OIdjeqE3uVEyvs+J9VOIRwf5n+kP4Gi0frwX9S+cRtWSd8ZXMRgR0tXQmMCu/YglQRzduQbgIs
fWqHLgvpSp39smqJ3CIe+2JbPhqUqF4BbzlgkuLvPaaY6xIk/tcO9PRCMY7ALKdBfMyZWdLMYdOB
Q0B0oX7Hjx8vNInzDOAR/njKUayA/wlv9wsWx7s7wLrSNnDDZXpuOh08/RPSfEhhGZeAB2Tcxxlm
nTxoqFTZtoRdAIFiFvaZkw1ZxG9bzKZCHXpolDKcg60B92DkwzMKy89L7/nLIntgtXF5sbpGemuJ
1Ix/Sc0cND8AIodFYjdnCsfzVNoJ7cIdMnjIqD0NkvRQi1/w97Fa7yBINTwZfbMfvuJBD8S742H+
furLG6UKYPzAtV4tcCMSvrpd9jZR2BT4tBLi+PeyyNId6o5QKEuyR7ACDuTyGMftbUnfqsxCxuvX
AUOJEN74NNbQa+yrUxYQgf3r+I5eiJSjlkrpzrOK5tF4UqDXTrmGrmhQY7P3F6OWlR5IObW8YpNr
UD/8EY//8y1D/tUUeqba7C5vzebP7JtBP6rXNEyHXuercnZGlT7nh4nlWqim/aBgPo61bHYxk9p2
pZC2sC72EBtEkKr4j/ggLBnwzVb3TYxM0uKp1BeLmHE9j+L2U28P35BcOl8JA9HbPEugOq1U3vbt
IYgaIyB9s80cZKIsT62VZ51SikcdVDfggGByrdOWKxW9ew8CfiJgxtwcZaVzZAEeU98WDGKTI7s2
6tKgfJ9ajjwA1YBQr1Y209cfrFCQfef4v8sskhlRBbMPUzV5o7Cjb71xIzTJXVkTDU7Mvq06fb4I
1z0Svn5qgjKZCWYmN5/NshuUo885vqIO65/B7YaiDzP4l2W7WJXcNuVp+tZszzS2L8f9D1WcWOmn
wlKbk4+eoQvy13/8bptZ2s5DkKh3i7byzkhDB2CwIzMaU2nqnrWgjBwSw8Id+eUWkyhzhQzBnTNS
jNH8YxXKU3KGk6KTSLSbM1CCyGLy33ZxUPhsT3DVfAfYmJ6gewiFhjuFit6UV5j72DJOjASgVQx1
jeBWvWySRXJUAxJckF1m9R2/DMecmwJLeZCLV+1qJx23CCmQpCSC6THfw4WbOXKr1WMABbGycAVz
i/MMkLakTwSGGeZuailT8+2PebdNNZ6NHkIo4ej02IDyPEi46dv3tZt1dTb1RGKO6vXlnZiuo7f5
DHprglQBLO4ayejwpRkUrwniSBrAx8laNO8qmmUnqbdPRRqodEoep9QGzsjvEzBHCEdGxH2jbENK
mR2b6M2VccOrnqdgIUdzDnYHXvh0WRSq4Cx7uvBfs42xw+XYq7uZyFeOw+BkebNLy75BN6sDOMy1
XLkZ9jOpDnkddw3qOkSl2r/MALbsY8yLYWmvnNDosQmVIYoKHhNpR9ETv/hpUD2VmQGau7hrLOku
CBb4sGcPZg6O3B+fJfJkWqlAmTCfG3SXnE99G9FC1Al3fQ+a8VqxrEypJKE1g1zuFFAXLOjuCR4/
vkDexAZsdkQTQl5HD1nIhnqoo1eJ7tRdFyBksilOcvQxwKcGyx18856ccvO+ZbrZ86RIv3g8S9Bn
zSOO2p+AWLjkoqEO2WKUN42r9eob7W6VXol6P1r3dL4Olmmx4WCgeXJCF7fLVjq7hQu4YWsiXrAZ
1yZSdjg+KlVmxImN4z7wPiv5njG89dKsQ2XRCsq8FKnsLB9RxCCwP4NiDTKsGJXumSYDMvZCTxqT
Y/eOfz5vtMvjk25ggNchrEWNYu4MxkuMFZAgjlGTJGLvs3U7BBacu+1QRttx5UTsV5PPmKvu4bWC
DwhPLlcXo0oS6H89C5DGb8pDlqmf4RZNjUR5h43SfEn/admm1N5mLduGA2OuW5ww1cG9LjbLzbcr
Sk3WnpqOWd8i9eIp56w/bBflaXtnA6I3Ib2vZj5gBjUNfFCLLZ9+RHsThd7VtSrpbX1By9smbSIp
uqjn7pmV2UwUaVVk6NtuKLkI5cZ3neWHdXBfDXxzCEybW85FT+QiavAotp6cG+QS0g5c+u5FvQg+
R7G6cecMPYFbRDVYzNH3Lm/M2aMOAAEsOyzCo0WRB7qwzDdpZrExKCxcB9PnXd3oxj2IaF8p60VX
7/er0XSJkDBgEB2zKSYDyyNQKimOH9cSEPhNyQFAXd68Mzv/uOPXDF81aJtvGK2GZmLz7isQi1sI
HJSdwW+4w5b0qeh+HN0A4P+7jbw6BYjCz6BQ3LiB8DpMoNeqTWwKT7ZYhkJvK3+bFoG6RYbNfvoo
HX1DtXGMfQORiV2JcsHY65Y/5ZTKtSItVVykdIEmcPiKqO0Z1MzhrIN3AdqLWQHf78SCRmije7uR
7fgdO/P8K7QDJklSGLB/6lRgMe4ClfcVM7M2zCre3EiavfalEHbbWl2uNamTvMiGa/+IPZPaaCpV
t9UfpnXtTVjt1xeCVQMYS111ftJUbe/7Nqb7Ge6KV2O8QKBN8OqPJmK0u/Mga2sn+Yk2TQT5x31L
KI9Gwq4nhcYNWHjQJHqa8G5UCq2NroEB+5hHvh0ckI4LmI/FygZ3kzw/hyNldk1d/Npt043Wx5yW
VvW1F2f32pCTi0vGU3U+nCuE1XjR/fye/ro03yJiXzfP4B7Bv5tKZfUv6r4fhLvb3VP+cqZqWpws
61uME0S48LJ9cXyqLdksiTMtWNW9IfmEw7JiRPLiREI5tF1MCn7rvuqft03benkZiTWp3gGoVXHB
aJ/Nu6aYS5RxbyXd+2fdvVQjbOFGtPswj/XqU0xGjBRDNgsUJswn6iXxV2gHu8yDnjqpVoGCi1jT
qdLsQUG/V14LR0DEs6OOuQmKJITlvZ1in4kqpg4GmH6UcGgvUt3ZC+JdcqnowcAl6fTyFknYV4Rm
W0/0YFfvI4dYqMffNOr9wAM1lbG4R7vYqBNgokbBcis04amSUx1JX8sjuZsv16afJQK9ZRDv5jUF
nlNSwxkja3B3PuiSYYs6vlrOw24qJVRmooWvwlmjZFfT7C7dHrrhh1sU639gpUomN+GI1nF4lQRk
NgZrwXY3JzLPYY+dtajBKSSLuAOyV1CMJ7LxZdFhqqfK7gamS2fN4eGveGmNGoI0XDH7mlGGVVkv
PQncAcaKXRdNtg6a/k2Yanxwz+OA+vR9BmozMCD4jC5TXSMxhQPVp0h0Bsmm5o6i0X5lYFgf3ADn
WqelkpfCdp9ta1SOxPwhrSSRnR/ofZbktmBYu7xzmXhH5aMGCqr/vz1Nw8uskiD2fErUotjYltgg
UHlvRyqFyqhwxy7/h9LjbARTxOMvNDx+dryIPIgiQK1X5qmL/Ks9UJsC1BGjTR+eZa+lJ2f2F8OK
Hp/tN9FsWEu6U5x3SVqh7qPDaUMWJyiLHEOf+1ZF2fGKVeyFFvsrplEX5k9AMlvYU6pbWqxqjwG6
83PGN0JGRsaKQxPOcSNTCOTipwEykFe5b7AeI7cfC0IIejDLvmHuH7NeQtTDqv/NDzXb/Sl1ehD4
pMutFrnmiBRjTytXrZ0a3t7lyY2UM24jOfPovv/g5bteogCTCSn/EOxZYfHnDA5u5xbpYCvQR9tK
nLvtpJOUqUnqlE707ZSHvH6buJ+Ehr74PDWP2Kq+FLb3NpjSA2kY6obKm783rYCNQkJqAOyenARn
jDMqLUCngdj65hKmzKrFZad7YDhYASonimcQzS6/rWUh12w9VC7gUOuwxtxLhV2UM5f2GjbYgNXl
XXoCP52Y4eScABd3hR0XXkENltH+OqwYgSaqwsqmR53jWIpcDL+A7mH99IpvzY/jjn6c505X2O8V
81ZrVJDQuws0NTMAtNS99uOADYtjyQWjDrHWfoEogsqmBB/L3CelTxMROjs57vVXt5zGts8MBfTg
GYWltfsC3da3nIFdV66nIpw2YfEXbLObjAQ7KtoKcLvkccczWaMFqSiiN/lX6PFEcjT3Fy0QGgb3
ukeIcyu2XhzRPYdYs1upJSCBX2kAjhT3lsG45n/dUFSO7Bcc0kWAudT+hRZpZ7E8XokQ3Hea+gWf
R3EMMkXFTAQqxRRqwdh6L3HXaCEGh9z0JJnso4Zbkail5AR64rCTKfMk+6BZ24NTKqn/7pB2ANcF
7kcNbuvY0btIjTWx3jgV9NvOd6Psj+uowUIk+ksXl4MHQ0Hud+fFu+YkfC2l80CusHRfNXO0lNZU
5TbZbksX0MpOoJOBEMtkaQ4LnbmHSn/5tMByVyKGd1HKdR/IgpNsD/Ohlj8MhRI5Xl+I+8pA8d+v
FI0Yhf/wmE0o4nuRHO09lnjSTn/+tTcapmG/nvZe0u/BKWNifUjesUodMzx3tkyaU0XSBoswSUbh
T/errB4lAraBXLIoq50JhUXGQkVHwx0iMz+uRi6e4RP6cFjNnEAZTPG8IxuvoThmz4Ejc2LIu7DA
9n5YPjgl7aOYpwqM8XextpWn7lLAZAbjO++tLXb1R7+tnZqqfK6JRFc+fof8DDoCXo3rJwYzRDLk
3Eb5cKjlKNMVp5H9JKv8evFc9GDJgAlSuMbp+kzavLjAPEuKNdOlnbvOg3Y2hEQHm2DqEmWMFrSH
puCfyyvy3CgVmrMBSoo9Vcy5bC1Gy+Vpju6kq2r27vK/4h6QTJ4Njtxq5SXDxFK7jnjUTwxPrTeC
FHQjH3JCSWcsyRD2/tqdzUIiiHhD9UE+zS7hg/BE49RF6gBppPvJ0V/8nGgBiio4qCna8pp4Cq91
gW7dYF3MdNyO2Kxqd40mhXWqO7+fakPqBQkbY2Vpi+a1B2gHlOXnhraQFPUjeKnHcpBQD7w9uyCy
WH0KLC3fpUMQdhPWQhvjzC2UkN0kFVXH27pKUwn8wamWNTW9TDHgvxLptYNEnKdTTpBL1qSyv72N
Jjun0DvBadqqdewzf1yJheUOTQ12PFMo0DNtn6aOeCZPWh+61I05WxuoWytuFgDSmxaFdgoEVMKf
GqQbJWXDeJ+zAGrkOXbSm1lfZVz8PK1t4Q57UFew/HL3dy9aEcLjXK8Q5kGuSb7/FGx+BA6Di1dW
Lps6ZTsY3SHlGjrpOkSnK6TmQImpMqDom/TAnFcTMTmyvdHwlD7xnUJ7A2OhDqVlY+I0C2wsCQpt
ZAhCTONUj32FQ4gtLCIUOHlgmn3D2+ObV8mmjUwIzubaG5UCRs8RNU940s/PKxQIk9cyssE/uCiS
Ohwi1aSsnFAknwWenAE9kjBxjMkzpqHiYzqhgGQyQkO6ayLk3oKLXC9uPXMEiwytePQ6OVoAWhU6
KnW+NHgBurRd6fkqxsCy7MEX1JCzNuSCPxtvTSyWyDYYn5w0DEn2PK1EGrA2xvgqt4oYgV2ePMsQ
BFbGc8q2/rD6v95mI/t/rjtlmnF7poOypjv3KU2tVGAgTpv+bjjU1o4y/ZIwyMwTaf9Uk7TbB0BL
ZKPyruhCcrZXDweoFaCcJpfsQoGi10A/bGkPazKGSslY1/Cib4EYIyFplrkxx4lt9GNew3fUP4aL
VVsJfaD4DEdd5OPMGrR2Mk7E+8Gop0QUe+JYEaVvv5wxYWxi7CCNB8kgNFPV5EUq6JEBEYet+/Z4
q1VOQ5mc30O/OeMBEFCwVmEhT4mtzQGF7iQXuLowlM4yt0vgtjcim6FLV1G0jdNKKf+02x80IsWs
4JyRvsjQNEjf6sKAhMAUp1J0So2Y6VvMekjchsOw5+P5PIj0jIV2KO20OYf/X0Y0InPsHOsgloYD
xKp1yNsIuybvN7FhakxeBUgLpDk4i10fol6dO4ADCyEQhpcMo5qZNS9HI6X1IqcfQFpmkME5L42J
+acT0NjVGqLOclIc06vxOFAPJzsXw/gcAP6EabLCEUG3Qpjoa4tegL9/0whxV5EX7Au4zmK719pA
rpshhjrA/oc9Us0x3n0feFU07ygnCxtr9WJlLa7636xHGRu2OFOkNDMv0nxUXvjn1S/5eTuXiOqB
jzP9oAU7fss/DL6jYyPrej4R9mS2FinPDWgvU9sjBQZVlSxOwsIoDnK30yqlGt9fNft5vM0kCfuL
g53ymZsPLzal9LRvMLnOzzW1plTWWlEeh4YvhmZliT1yiZNBN1o/9ZH4gSbzjA150EyZtx9et9U3
L9Ft7rywkxkQuIxahjVT3BgjNXc/2bhN2BHX5S9tSZClBGrpQkXHBkENWnpp+UVWAteJE8gVfkTT
XTBlliw9QWyh+Tnkdtr+H+9GJPDADA9HWBgNWquMJZvhf9j4RSG5onTOxYLwnvDiDYAQUN4iu8az
uXzV6E/SJmb+4McSiSa6Yva0cp8pPDTZunU89V5lYFp23J0z+h6RLqaC+MTN78Jwy5rWeWER8vMc
37JAg3o4rtxOeWjUIF3iUpkJfkD7yZ1OJnmAXzEeRT1aMAMiOi5tF5Z28FfYLWnpV/f/DcGjw80S
9aYlAduGpyaTawi5bPoRIDYBdonhqw5003dFDTYtaRWzlwuRRtLGQyqTu30bOKoh4pEv+XIsDDcC
PZpIeW3jV65ytRieNz4nMvkm3bThRLuIVocnI4RhrSid9DzjdHu84k2xhMHJJk+F3lbzEI9Jjo5o
rmMgaxlFi7RCMGCtJuQjFcIAyjzBNeozoC2SU0xMZgAgjt8lkgpELsHV4qOjWcaCG3gZJn5I/7JT
vAbg1jGCxF4IpxyGLiWIJRzjVanPxPwb9x/RsU7hrvvP1dCPDBnFu3pDxUDUg4in0AwtyvnxQx5Z
qFCc4rPx+JSJSEHaJbS6xNwSbVHfaKW9Xixv3KxojqJWBivxBAoGrvEVgqNhUQAqqEp5FCa8CkJ6
ZEuMIHxiSAXa4F4ZQzyOda3R+/RpzS8ZccD6Q50U2TOkXGfMnW9W0a0v6bB41rVX+T1n22363bw7
ujYm+SZ8Pbccoldwy0Gs/sww1M+7z1w5KAvUQ7RTjW1l6fq3ZhCmIXrXi3gF3TMgLpPSp806MTC9
bNj8tIG/+eouqHhh30iz/LtORgyABBWXPdtiWadk3WXHdSJa6k7wi2W0i+lSQV8TDovUs7cF1noV
Nwal+EdYw3JwubibvhpZ0t7VAroe2/DtAlwORGtgzJD5csHbFNO5VXXpcfGrVrmHEFIyUMI4XKUW
Q6Ot8Xin9mYO3/Z5URDYorRGwhMHvD5msl4kQBvw406zP4Mo0xSG6zDw5N/oNJY/JZKlaAZUI3zp
CqWjQH87BOOCpyxt0b5e64/nZOy3cArJPDvF7UDqSDDjafTzxBjnNrH3nBqGmZPamfnSZ6u5aqeY
71VgGpvHi0f1pPh7u+tnTtPFdL83IzQbLufm21YE0Fvj4YrrG+I3hpqadeyQZ+L87Er+5Us5H79w
t+yP5RTXfsMHjsJtKmpV+kg1f4ZszDgt+pa7yyZmmD2B6N3IUBCseQ+iX8+rbGrZ/lYw9gfVJql/
Akdo2FXr3hD4YGVYj4+ds3ZWjgsSEK+S1jLOJRxmc9p1lVCvlM7yvX+jxhoFGvefABX+u9oEdP39
GB2y/k8WMPUEI0JIFzfNVK3qMwEP1hx9D84fLf8LGFZS0clg/NgYQqKJeQwle1lzShM/GMhKwIy4
YoVzEeG4TVuj8wVWfw8r+BtFW0a8RtjBS1m6cdMbk0mw3MEQKjjVtVqFL+i42iOUSmxN3sy2rQQ/
Bg33Cgwb9dIhTemU0Hdq411kjMoOqaMWXRcYKX0GUPUkoC+Zs6uFfIg8r3Evv93+lNswvP3Znbu7
rZ6VyT8zjUhnbkLopPAI9GTYXw4iOqtfdW3sYmUsOQf2jdM/O1Y9whCrJxcJDca4NYp9sqYiN5Dz
OpiV2M+C4JYBKbVZ51EPwCQ2vQUWsaIw8oknZrnmXtksVqBZNnRmPfdZqPyYWsa7m0C1oDcKQrG4
pjYmYgJbuuf48ijbNj4MlNXIR9M48J4+4VYjSfMVkH6FqqYCboegqTPcL4P61P198owHyyXE90FT
+BpIQhJiwqwsd5wNa6mS6j+WtpoSHazggspZPmMchx52NUxo3mvJJSX0CtiHyAw2qyeBaYG/kd8U
338Sjiy7wpFP040c3uVJCwoku86z7cXchCSI1bHERBPBBH2o0kP2ZnjSdjv0oxGAcdt8cLJ5ETVT
ezN/FeEMR0Iivsn1/yOnpO6Xb0+W+4furXTvuSmMisEgWJaVLXF+wGZ/n6OkZ09oB7bo05NYJCt8
3FzAW78yGaBFIudFTDJyLAJD2xNDTbZJ73FRzjHv4sgunlOWZarW3lGB1euegFocU2qQvixzPk8g
Cbs771F3206Ga93/e9qi1dOt6QBfwE5feXm/V2eVfg+FjZo8MEKDEuw9rzj2xYx5D9iqKqM6e2uD
5UspMijl5A5g5rG7s2iAPOH9j4f0jdGXmHYA9jmvlLuyia3mSDTlNhLcjHFFLE0GwBCuK8Aa9YdL
bLZ+1eaJQwdr6OUeA+49+vmu0ctdL5gyn7BVdO7mtpoXoRc8KFj9DObGxIW+SydMziPQP56fWHFp
KJ8rzxTIVWK/BTeRRb2rGOT05UJZ3PxLybdXCBJMRYA4m8QQr1yY6eHG4UTpQ0J2WwFQqCWZ8z+u
LMejWVL3K9Pg/DfPhFW38qCUSnH+wzL6PB0Hzf0m7nKszOY05gshIOaDBw0Uo2zbecCjAnY439sf
BCNsygrZYScfeCBH+/kq2qGnHKO/wKvBmhZEo1hJHjNmei5aiwHJxGEYP/ygLJ1gUnWFHhH/BP8q
e3KGqsQ13DX9dRl86azk+IH1CZ9GHtCXjnI5KWduFhWWAafEhKGos58vveSiTd99MlRknCDUTqN7
F6HLgI3Yi5iiM8MngwTn2thaa45B5gBoxZP1+5J/9KhNwEvCxdbSfARpAzguwc6sfTLTZ/CthcCS
S8HtWrSdeqhFHceewpXIl8kyf4COJEiAoVOl/Ye7WLY3xCFvE1n9K1HX9YXoCbMb/K3Nh2N0wpLN
JNwGUupm3Za9+DND0WmgFLKD2FvXdMKHeS3AhvpsTXOicI0tCJXjA4HTfdBwINLhdhCVbveyG+WK
wLtGbvNs15yY0cRD8Qstu8v0weCRskmCcvrpuinJFlyRXxvUOcqhxSABH5qdIwR2Dk74A77ffBZU
pl1uHD9JHbGXbLXeKZsaLWKI+Zw7Uo1xG5uXWYDo8hbE1abQT9xYX5p7hCKgwM3aPUGwENiJX6HV
7p39bYn69mVpQbCEEGTxFIDAbze+mEfafkzXzhRDJp5mISJDv4RVgJF+O2HJQQEE9Y1rPlJGAcSS
C8g/J8cDeoSnucjVdDWDqddHr/Ljx7CveF+pcptFW9gXoySsakqwxR7+auDW5S4zUBHb+j4/nlBv
ht/9Yvp440fj2C25H+kecgmbl6Mawqt3XK9U7kcHeKOe6U9z5GBEBCSXY7S5K2UFIL8goG90+pQi
OOMPhP1nIKA6vyQP6UofEbk1UTKoL3RU6ipMYuuLR3+XqUVVH2R15m3wPJ8MsNCmHak13EsXowp6
HvBHehAfRo8d0K4M2G8jomy9pI/961CYHzPmv+XiH17Jq8rg30wMFJWu5rAEosktY8M2tLdEU6PP
hGM8b++escXfNillAY7v7ZMVQ9u5rjeVI1JlPAnn6boZRssEhRFBxa7+ZPZKSRAZyLTZc3uOxuzH
yinN0tlJc2OWbVfZ5ZitJkVNAUF0k4tXJJabeiI+WCdryUFPBfTpTYbdKK+ceqaZtIwqeYIDR1x+
DKfNxpJRjaONt3zMfh1RoAdx67zgs9q9B2t5suvrKIH/JoRuN7nrjmG2F36+ivLEfME9kyOhW2No
udFSADe451JyLyZ5uuqRP/rhtTX/Fnt/EW302TkhyA2HOCIikp8385FVscRd1VEkTE+Ueslw+nvS
jMx8Qzw7ACfwNOXbFaSr5+3JwhxSwB6aMpHOmt7BbMYnhxVxJc2j8ih3LAbScOTxOmhqGSfwtig/
AmFnnHVD7yddirTuNwPfdcjZD+F8olaeODA9L/rpqkIx4XGqf1k5K3X10E35jqYFTpMH0bsYNs3T
kN8/98F0cIYV1xozH1jNUB0QLOH/MTdsptoFfDwlGWbFPTs1NwP/zgtSXmRUJI0y4PBQ2RuMEMDd
3GXUpSqXJAhAAPj7I5tYoGYgzof+Be91fMlaaN2bGjieuddtnkbqBGnwKPb+4VwYQ61YG+9l/Y31
zOy31WP5/3fFl5BvQRs8sOQbhmONVVBVSOIMhTHJa85hZU3JsTZG4ADzkm/xH9Gnrc6KRwhNOowR
p6AG0cIRfZDd42jIeL8inTuSsGAWNd7vq0Io8z9l92mLzGLUVQI2ftdfiS/ddkiroKZRDZIfCcH1
gv6P/PGaKtkvPHmP48hjOdXm5dajEBz9Mt5FYeiCvdOuLVmS/1MkuRiASTuN/xsiESeqxhxiK3Az
cMkMgXKI2gd1zZtlEFHTUEpcSHAl/6HBu8S0SlkDIZGedXdeDPemrVU0zUf7yFSUGmrY+5oWfqb+
N6Z7sTay+Q1c6KZUc4HZUpydRHoK25LwLQrXR1OhGGmHBiimUGneDEIn024Xrc+b/XEv5MkKYgqw
eoyKNYb7kQpZ3hYVMh3SrVdzupI3thnAJpkvPvUVxOlWUFPLj79E8XspqOZ0lZg7VSNbD4owa0m9
aMeMeY3n+pfugb7J9S0o+qQXgPqCSxBF5crf/SDzwtGEPcjAA39RmQXEBnrzPlQDTXmsnJ2QtIp1
h+23II7XLpRK55T8GPH9WZ8wSzG9TrpfcHwAHEUnTy5bY9EcYD2SbTUVNTJRCaUFRDh/S/2Zk3XQ
njN8dTJbzVQeI1zsTAxpB95eTJgWGCPLNvQcE6Piy+wCg7SdeHmCSgdg8QmARc5MnujrzFPF3HSq
//Ck1n1JP8lDbRZNJqzO0gxvNjTQBzZvzpSnlrQVndpfjEHB+32VqngzjVXU+thq9VHIV19bA8iX
7fjYJ71KtdftRZaw5HRMVJRZqs6PFxPvbRQFzIDdw4i8hIGp5DZ38poO/UYw8c6V/4/Yn4gkq0bl
xTqlUZ2NP1GxcF0Zqn3dvMYB7eocuaoqIMk7lh/N1JzNAKiw6l5rH3dyJIagSx+LfpYHoPq6itqR
3AZ709zygT5MqAvrODv/gbrdh3d4ou4Es5ViM2ZXWp1v5HFq55OH+EIEk7FcMNrWTpo5uUavB9GU
b0yU6srOmDLAydu7jNydUQhz/6iSksMoXR8o5kuv2vQ+B6YeBbubCYq1wQvvY6GuKSVujP0JuqJc
nrgOtloTlPlEhnRs3YWR6imN2kJ1pF8gqmPzMKBUDIU3oHdZcZgDkvrddgP2IhEjEK9pohLKTX9P
4NDglL8Mf5ObvTtvuauHfDSsJBZCs8Qc3be5WzfOXFEuUhS5raLyw6XhVGHqAg+k7XeWzg7X8V7O
linHbu8VnqE9b38CDda9/ysFbZ3jZalAGf7EQwUYJqiyvJjV2OMwgbQbRQLC8Fi2RrulqZEmiWZa
59BKhtag6hB873mdEEs1bK2d1Heowv5VSTDLefUCxgFg1R/HYiWqyqaIySPc4SxABIN60aoxUK6R
a9UfmFyLQS6qU0erI66EvvLLFjym/J2EMGrzbNAo+yygG601WxIy4x9n7pgvC6N3bTM0n+wtX6Yz
mFwNTeK/oVUBWdppFpIc5mCuyMOnMUVG81SkEAXcmR/hZYONamgHELbQdEKCcXsy/ueD2C+4wA5W
SGWTr2F9aIJQY6tTkfTLb0EQJZZsRANTrTAWCW5DuFDnJIGFMy8D9VICh8twyh4vQeQ/M2DC06ID
w0VkfSubwbVYW1BwmbEFJjp7CGWAkQhEwkdqmi4mWo0UN0p8hnx9FFSw7S1RbdMUO9h5JcRjotBk
8JJOhiGFMUNXi5NEkTymasGLWhbrEY3DnmcLVHhPmAprXL7/UWl2b0IlzoJds4aYfaDYfBQpHx3T
lgqC9Kv0utnY3hl4AYq12mYlWSi5E6+GHQiuUWaqPyqFOHac7Z+GtUdS7Kr1SpF2n0T1gsHNgYna
NBnyOjqwHM2BVoOmYXPd1buoR3hxKUpuO2q9s8AoG24EKf3M5F4oOcUrKG8mK9SLVjuVMs3y0SNr
c5Lq2bsMvHabZ+lUzO7rlt/YdZ+UboXg/yUm3AGwn/DdOReD1VA8jtwErgLkJHzvK/QYh/H617qB
Xjv6SBy5ysvrkRlJFvIOdk05mrLuvLu1K8W5RLhs9z7Pqt45Tms1rzZ0j7i0E4UqqqcFZGUkKQ/H
ERevIIoKrH3/39wT2pYkEWqVEMehU94FhRgQITkx23IG0TyNXFZ7HElS668yMwZ2PYQTklkAevAg
dfxRT2+aRn1jfQwyLRpWhU4yNtwAFmrcahVx8aOrPmmN9TK/bP+N9Vdc4d7x1GNh2bHZreWraEWu
kZ6AZfwOawgyshcYGSEcqs7fhPgoiykaIEwIdybQiC0f/hcJXzibeRjRjaUxvJyPKFLQqe1v8LeO
1iZAs7FvhJsnF8gd+LyjiNuM/Py0MlSR6Sr7GI3QXVm2Rs/HOzSX2ecldthUSBbEMaTF9zMJb88V
EPlxNDR4dfjLyDdRSOHS0MQb17CcCtmnRFSnXsUKa2gy52H6qsO5TWwnmEccPLjcTr/gX92Srrwb
YB/L5oHcp30UUeOic/ACm9yqmYaoDYcZtryBooy27XWY+IV24aJov2XdKVzNkKtgLaImFf6/pSyB
9ePDQEFW4NaXXtgZm7mh2UNrdeeypmQWppnu8hxD+zHNoq14CuduH5X3xMbjPbPj0AHmcc4TnSfu
ePaLcsMyXvbG00TmSqv0Eia8Lti07l0yCSDlJ01gfOAaYws7rAlX+KrpCaXBGWeG0Ty0/bB/TzVG
QZaotlJcSbRCsKZclpzDbblYjisc0Uc1GlfEAdQNDTrwMnslydMxg/8VxQuX9TVUTZ9kbzSZKkrr
N1/aG53a4JzwNND0LHmscG6Gg3S/kssbpqZYY94TfJ6h4oLHn8a8fAFavzD4sOSuJwZUYhjm8fB1
kVnHYPWTmiffcKCLRfJ+0AaQJMbtEV0hJwgrWQh5R+xz/aQpDkZ1rv+y3Fl0YnxJWHem7tgey/B0
3E4MSLOlswesM8bC35v6OFo5e7C6xRSsaR9OicI+UWP6/o9MVarGhy0CVyfEyZ4vW/fgs8/t4T+C
6cPrJ4h9n27dafUed5I/9B+CTdga0k70K9naJ7MnrUzskUGYlJSQGZ0/Mc1wXIZpI9ipJeQNpsUK
zsvQt9aCWPY/OOxMZERp1IolCmda87Y/XB5dJMMy8s7Hu5nVBh4lIRvH1laLad9EtzTSADWTJbuJ
dcYV5lxbI34LysIWWITaT8fV2/3WEOQSIOw8NsgZgstmSn3un1Q+rXWdMKOMDPfdTWWMF7rQRZpb
RdCGZb2mgCgvHLZGi3/F5gIluPvqeKUce6n4ydrQYA29QqalDURRjHqHV/kjtT+Yao6nmpfkutsi
/g07c174C699rY2PDUiIvOv5QAybpjFU6RqLJHRwv9V+IZLXG9hriGXa5YQcn4mcMoePgfBlT7wS
bZ92hs3+Jrqr51gQ/HXB4zULgCXFuOQg+tu4sWMEjUCd3pjRzcgPFdae4owlL80CoxK0w8/eFK/A
6+rnR7lSq74zQwumjNP1a2MQrGx/PIQ/8AwKUsSyrt+hT7Gie0lj2gDqckD81YVNZOqCRR+MeDsK
+WEgnYLHX9d5Dk2OiWO0LJd+DYom56YPYOq1mEWsSS36p5aCOFGEMwmBSmtk453fy+h4q13jEKga
wXdyUI24CAaTEEB5Q9BLtxCIXGyf+dn/e4A4lMwrgGfF7eYf+rl0qpy9lyHbRtR9k7T1dAFq43dt
iCy74C/t3gTzp4JX0jRurWtjDMVm7Q2be37ZL21ftpWzgh0hhXiCDl16yXUfNDPinth10CqxLpIK
SUAaeccrLL+fUiHMvCFCvYmcme6lGR5WuWwDp5lhXnrcgBDxZeNKNxBAmSltJtdNhs58UvuNy8du
iXGBxXID8Pa2n73k+/RUeso5BYohK3sKDCFWFKCjTel3Mub243McsR5sp6GL+ZhNXfMbgbO5jf4O
wIqNZ8AjsXEo6ZlfsnRx5UPuIYj+gaTnN4rzWs6gwqdAn/YXjR6WcEGA3XWAe8ugSoITscl/z8fI
NbiqjBxpaHrstHi2OcVvgHNWn7Kofk0jDanqFzBRPaMhXCJSUew+quP+Vvsiec1e6m/fYwSNq5t1
Wsn8Qnxnjd/KM9iviREPkN0G7qGcPJXu+wQxyi2+LqycXFD7K4J4YaOTHU5DvIhqctHk7qsbDkum
infksflcw5ltEXOnK0LhGjONbaHQTA3/VMCTK8cFgEYNDqDxOu1VpwV1IvAF96EUGzKoiBRSuo9e
FzjESZ2/oIUJPIuqfnZkBiDJmvve9abTFivUIwPmZD4ETnhmolZNpcxYdGVXT13mbYESR+POJgqQ
oOUYrhNetuI9S+SDJoea2jfbVmEsdnyLC6x/bUgpCiLK73esU47nmMskxqnWzRgeewm0no9GKcQ7
lW5XD50/VGn62icdoFu2GliAiRnpD56RqgpSVv3aWSyMelc2BHdq9V91fDkwlZdIGXQtGwuwevHh
JuqvNLz2xaw9Nv8ijzrBAe/DRvMdwc+k/4YCt6uwjvfa79Bq/uLVgIQtgi01RbJXHz7BDOLtyko7
quP/v5pWssI4d7URfd6T/FXM8t8G37ey43TnvGRC2xVqsGlCmgr14MaisEaOsG07Ean5Iad8B9S/
GNhTcLPFgTLXZvbjI+/wpd4pYfP0Tk/TNSh/pP5Dn1yNjbNXLegY7k9ascb8GxJUPCNuVRo/wW2r
k+X/Y/gcA7JwQ3ErC8YJbk5j7j6cEhUm2XaOrgcBjHB47i2T48DGEGqq3AeDiSaVMXtcxRsTuXJ5
xhv6pyDvMaQBW7bs/qASDPQRGMCY4r8OrYr/PSACR/YHgSMZW9A53MA9fBEfA3GoDePg1t+fXRPb
WVRggO+yG1VYPB9gx9vwn53KP7POpZq5jNUItxBCOBJpdxyD02Rd18NT5LBHwQMPBal9/SFweN7N
quhq0nHpHWC3KPRItw5hv12f60iJhSq+RT4hHh2ZTwIpsTObCcc/yzfNYJk9VhqmV54BMlK3EUTa
6dAGznz1qyksl+owm60Vw1XSim3oABqsuGvjzSsRJaaZvwhq+uNSTR7WwK6wpT2SmRvpH0MLXMLE
9KOYe2sResBXcPrq74O/+6z7yzLfK0ooLX39oSIOVhEgpSlHBxfLdFE52id06qKh6/1i31Xn8kBu
kIGoXPB37dRS08F5YaDI24pGkxz4Fc/ROQli51sR3AhyhvAlP2Bxoltpb4My6cuIFqzmzf/SThlQ
ndkg/j3Gw/n8AOioWOG+qNRVrVdJHPGbZjrESWG48rT8KVO4ZLschTtIkyrQiJagP5RmRkZOf0oL
FBopNqi12GgHksneKu4Yadl0QMHI+AF4BKXGM0mX1s4Nr5Fgqoiq+Bpj91fyd7j8+IkbWxz/Rgpi
YtuEwTb1YaTcT5oMpLCYMtud40vTMZ/srKlOA0Ef82HA73JXqYXwdADZNAhiHLJNfM3DL5fOe96g
S9/Iyyft2VDvP1W1I8MqO0vD+B0P9Cuh6C8TB7qitlPMg0HFa7VM3CFipRxiixf6hEk6m404ds10
o967xd8YVPYNDva67ZHDh2hnLnYUEq/MUSgisTOAPUelc9LIE7ACtk2UcJYqYXGwMiTTDXrpg4L1
2C5hRfRolrQVS6sdYQjEuONFItJhp3u/qeasQy48hwU0eOc40ejllqhsImVKUOw43IlWeT5dZnQD
2KvsLtwpD/rN+SyJwIAS1FCeFHJnmQNyLp54TLGDkupSeCvGKsNgDTy2a9xMWe7sh63qKGGzvZ5A
10koytHmq/qn/pKGY0aPgJQ+6ak16P7EMSqzKQ1siOi3ml8WDF3mmPXqZw7toJec1d4RVtd1IyRj
oCRkxdINa1PM8IPSCKazWaDQ1HQiqQC6/gXhgS12BfYlod4DJly1zhQEcdwJnSmiTqgX7RVzwx0w
T02pJ5zDI3vT0jluZeH5THPDWuNQaMXVRDw0JrSNI7zr1ZgOKsLXR45qEhcmdHY1dyrGeJ5DtwJF
e/66mwArrFJdVfyUYR8aOaZ/kicCPz9khnLrSBUfwGSXugpjFIBi1cWeKba2X28q90SSmcIi7VWX
pdgqC4hqFDkSAsBvuaD6k06/zw6r265vl8qnXfVtb163S0jhNNeeDb8ZZuvXzrCf8h0vihAJuWYn
vKVKQGS4YL27WA12hVizAdmmFdCPm1KHHW2AhqmNMZ1hKFnWntC4AZmHPaWPMzhc9xsUXBG1vr8C
vmTCOMH8Y3aSXi35bUjVtPzIZcvdidtPfe+u5Ppy1xt0HV4mUH7o/8vb6xqgKgzVZHmbBuZ7oByY
h4dsApbAe5d/F5VCR7Qn09WAyLGwi8q/8Nz9Vw+6S3ygloFXPxnSCwzpYqX/AiLNUVRJQp5TEuef
PZegOXSEXcCtrXTtgTpiyYvpnuYylT/BCn7mvAZsCiS4H2bp1xw3uzOyJW+Tm4I1ZG5Uj3LMq75a
vio1BtdvUytsw0+Bz3f5Df9qWs3X8ClwgVZV4r8q8P6HBZuB7+dswH4S5/o/f5lgk4dCzEC3ftzd
2xxm8uUMX8jYzgdEvBPxQqBuBur+nQeEXy0Lthwt+VKKai8V1rOIzp4JSxlSvvmpWr3DS0u8htOU
ocXImKZ4wBpKHVg/ZnTftpCg5EYWZcrXkUyCIF6NcnfYwqfnS7zCKyrJ5mPBH54rbphYcCOcAw+D
6STT5qHk+WZYMP1Z/hmb2j4BBv5d2bDTYxthN2Elrx3/nKjK9UEu5qpw+LmybhBozevqFbzy63pd
ZyVihYdBOfIgMPDcZd8HvKH0SwjqSjdWwLFk43uKudVLQGbDRD3tI7RoDirf52rwg2HAkJ/0qtOi
fS9Fmap+bJawxTHIrcse/Eqd4Gz0TOCMWXTMHsv6Z+kEgDL168RuP86ekHzDCgPFXw3Frb09vDf0
DIikacTWFsPqtDyw8/iL/mjOZJpMk7ZBpVIMDxJIx3ZUeiOKHSIPiDFTyihumN7TlM32ULAPWz9e
PBwnM4uXONLlucQACqPlL+J+3+ZQQtiy4AmhSxejMaBH+qO+Eag2rBPzeKaXfv33CXVY/xMxkE+2
GemRerr4+DsTIcTjpgYkuTJumlt7htvo+4+L5IYDacaa0VywqJuB54mM23Kc3PO5rVomPMejNCiM
VIBH3BMFuh38fi695WAZ70g+lQ+jgtWyNBWVzdb21NUV2wkw5XzszZb1Frl1jyNacpsNWznUmvFx
S4zXSjehbrT1WaDCKF6P9l2dUET5xG1mfCw4TDdww/kJtTh6ICy+efBkTMqRQxslVR8uJp7l5khP
Pck60lWu9T5kb7+7AGYRR2b0tcM+tHIPTW6Clw/+ZyUhmcAk2wth0VFQ56TMh1aZoU1u0kvetpaC
kZd13jndavlP1ExpgSrwpObccf5wmV6/vq+wnCKFkHtqCq5hCdPncdm64THcETWLG0MZXqMbrC8W
WlI2OQlcBYQn2mvMii5DkVytesdq0CF+fL9DjuPzI/4GitAndbKd2UkvVoLBrvaV7o3dJj2sJ7mc
2QsYTL92HEG8bnPRbavupHz71yOj43Do9M28DkzRuB3bUAf23PaSJwLCXEZ0rAwDyWQhXJOn1ae0
ClNKRY4h9uaA7NSbrnFWc1nuRHWAQ2IStb4QX6AspIxyzvIAXKdQHh3LgooRDusTJs4q5IChy1K2
XEbUKqujERN5dLAGKtvPWZejZS2bq8hayUnunLDlix/W1pU72u2xvEFDEjGo3rDsv1s3yB7ogzx6
XIoA+BOKjm/2x0VTZCH4qBQBLDg3pP8sL0zCdMy8TijjfWZN9xmS9zvrlllHzO3nuGpyI+XB78gp
yTCkxXxd11mgficUeLRvjavi6Ng7ie4oI+gWqInk5h5UDYhiM4v2aniKOgH+Cmpv5tgBLPUWUO/j
reOql3rj08Vs3pofWDaJjm0hzAlYNc8GXAam0ko+qWhkguU3JpybseA3mO7X3stGmxr/9Ur8ixPR
vYEZ4fqFuBHS/06bIOvNAVR8By5msdozts2X6vS7FAy26xofBAObcn4OyF/NNG4cxiQRmpqBexxp
BCPsBccpYAsSKX8PMhsZbISjSWqBGKGw23E1bjY1//224DTsXeOwI/1XJTiZwwyNTY8mwKLXlq1C
lHVTOnfW0wQNz6R5ah27k9BIRrOwMYVVxQflUlrGsclD4D4dbfoVAR7PjIXYq9acAgvv86TgYod3
aTKL7d3BBOocgkmknvTs2wWznSc4WF/Gsscoa5lg4kFbh7amb8zZcgIxXj4+OVUcqg6MSVep/ypj
5kdR0fEXwCcETfZPAwuJpnYWXiCZuDnCoFqIHXq05hS9yR73sQ7IsPe/IW0yph16bCUU3TX6ZrJ4
UZhSwwGfQtSiakYZO4e/mfQpKN2EbufRFrQe6g7bWH7oeNlMOttXlL3spYxQ80i2IzzBasNv7Mxy
HQIPAm5CJwbjvS1T9zVb62deZMNHq19xqT6ILEWzVNixzz7hDAEDcWN8KAYQu3FmzlhI+SnPiNE9
PqcDQkER9KvmhbLuiUA3VDvuSxnASZx2xcRMYaEhH8ipnFXtX/YSHZU3Q7KslVY7m3vBPUbZ7jET
ke52rTteFhiHcHfjFifDsZI2H32nLPu8nmkJv6TtWUerPzZ/rAUEg5QJ5x/qadDw+SKxvORATCGc
1ZMnpkmvHoEuiNjkgKnUp8v0/Yq7l0n1T2cO/dQ2dnT6Qp+ecZG4/BRA2b3GF0XAobKeGATmL2EI
dJvVMDnUNBX7ZFE3JmbiOy+Ce0sps5rg5zgohI8qhPo78l+E73ks7TgHuSgdMP83lmefe6latNvV
ZITrDF0KJ0uXCcP+4J6L+YyZgu1h+bDNqAxoI9hOCapAgji+bo0C2QPnluF8HoWf3l2Mun3Ouw7C
XlVQPZG3B855e8AJRTWplvBMh/7g3+aF/5GUsRgBlBsQ7oPBlsOjasM8c+gmcYYSPObsxSEtPJao
6sgRaiOmgBupf3xwXnKba4uj9gh/KlCYo0NdFU43fLY8wTFPInEEs0cvJsuM865+DuwzsfSlRVHJ
5lLEElVdfHzYEg8Euar+zD6nN5+dd6Jsa4wvxAdxQiH3pkZeZQ03h7TX2jzq+yGPJLxtAeWJ7Nv5
ZQfLwmaXfdiCu3eRl1bGxEZEfzB0Hk3LpkYevu+C8n3r6Gtpy/EiDMdcs8KD1einqb/6KLnTEG4d
pZwPWTWssk1bh4AEHpTkuOIECftt0Y1LYCxEsPSzSz1Jn2OF96jeJaXZDzIwq0JHEmUnggi7ycpx
EC7INiA8JxWCMTzZJ1K5xgE21hXycLHaQNd/LSC6m6JF4XArs6VjikOIwCvDd8V1n0ARBN61maWl
1LPoxzzEZwKk799tWe348Uy3Zh1GJvf/QB1sqD8932Qmo3phuNY5OfR7XVnl0c/o8hb4dZNugtl/
FbtT0mtdLs8OBBvWvlO60dhSTkEEsnXkrqhMmjA2caqWr687zZp0LDqAQK5wUY/GU5feLwdPiSFF
PuYIYv+QVJQwZXUc7FVFj7VpHFV2vZJqse4Zr27iSYzMmMmN1+f+xLYlA1Qkdv/Xffwg6BjTXDqW
boFkj9zEdK9ZScuYiQPqcFGb041vsAvr2KTBMpy2ceGAtzELc1oKORpXLx9gYfa/5LuWko/r2CNI
FfUG9h7w7ebFlQm8fmvr++YFH42Db0rcH74bjtrfH1naGGH8cgdFiejLjOfqu55xQeIrsWbFpLIe
SeA5Qd5y33kEcnXwIkIwE8/oIy/909F4yqRpjjmIJBFiteJVJQlEsk8q3RmE+qSr5xigwOAeXWPR
lGdO3oYJP+L+p3RC5hR1nMdtNIl3WcBJMGg+2lpopiLYjS4McGuE9SNYwADAxsOtSa+oAqZr1hpO
3ReeaKifdZ8IngTTGd6Rn/vn4lIMiCZd8r6aA1JoIvjbsHedqT2SayN7TuiEecCnMe0m+PqPRVUy
7+MbjfDjKdPTKpTSFpop5FTluqOi3P94MlrEPq/GRpcB2A4ftyCx4HlYM5wrW/BBy1NwhGPZiNh8
o4NxOG3aNETqYu390VwqNd7WQSDgYMJvfz8gupg9uLM4eIcIDxNHDCaCpVjXqUqv3dk5Z0Ks3PBR
KT6dopUn8LuYFVhfhuJkim8WOYegSpimO3XIEb/mxA8BYixXWZB9P6h9dP+A/xCCUqmv9b/mv/Kl
bYvzvsa3jBo3H+vWHKEb+PyHAzFELo2aNKRUZomMYjZI45wyIvRyhQUg+RPda1SiWlXP9ctQKrnw
LyDLInaeowkkt1CwFA+/PQAbV91OzCbCxzV85xpW5b7cRJJhMrK//mTlIiSeLrDwNjhbwnAD88U7
/c0QjOp16Bjo7f68sWei/JpFK3/hdg6sD9sjjd6N0qJc37paygyuKI8shXvrAbtv9LfuiWkTmmj+
coLoKPxXxFyfABUi0Ghu3J2HbN7WAHjxjxHiFEZNZCTfsmGhE2cGgqhUAAO04ewfY+PZALxAsfVD
08YVhJr8Sb2GbxIHwDp77LhdVcQWCYpcy6G7KpfTlD2X0L5CPWGDwaRmJfk9WTwqtFMLUZ8Nwbs5
v1ArAW/spveFHj1MNSQ6PnLBAI/6GxTJWTgpb6yP/27Y/5l2fUxTteuYqIcRoVLoI6OsC8wiDfj5
XcMvSkr+Z65i1JSoQ+8/y/ZHNBey8bC4jyD9LN3XEVTNYiKZ/05fSqjp+RC+SP+G2W3psNkPgJVX
2quFLKJoAf6YqBjMvBWfrOcN9QVQGfpddifdWbmLM4QbyJq7sf8PJJYQLlCI1lRmwgQXzYxulUz+
/67mldrtSMwrxK0WZitVX6Dfs0gRb+io2c7EVA47s1PmBguFPJnuHiubw5cBJiGbSW6mdhcuqDpH
CdLzhtQO2fjXoi4N/cuMLf/7dC9nKHeJspiMot+PKFzVqJXI1j24z8JAnOPwhcdb+DBUM/gZTOjc
Id6148Om+7T2o2hhzeszuRQgbHzJB70rnsN03049hnWYVDT5BRiVTjv5scam8/0SVfQgun5YEL9n
ng+bpBWECGWdJJYOf9ElPnrjbOVfKG+9MNdaRTiDjVYo97NESoLI+4NE0zA0QSURj/LCG1AZeiUI
cLcmDOHe/iV6EembqvrVMwNNARO/UoKjHMtxsxuQWc0jF+KS4yDYpsh5N5xr+TBXtkxmoFMzG0vg
GiyEUWCLUU/7/Yd7jW6ykRu3zNheeDDWlG/OMIpGl4kzBkNEA6D/iEbgWSM4Raop/69KbXHQxeMk
nc32khoV/Zb0PkmEsCFHUDwg+RrW23AQi5YIFS6vkANOB5uCCcgXcnBq7MSJnBxlJTe07NZjiokB
9AlQguTKyUqZl15P364rtYpNByf3sNqV7rYIDIRmRRgjKJb6zZv/TkcWP7xKvNtehzyL9tDRRreL
JWp+W5OHFes71pj/k3vKD1oF+ufbaufYlJ8T8z5Ir7JhUA3jD9fFKBkZEEQpxRry7tDcd6BCCPP/
FZR8bqfSO+wRSaeDqjyEKp0sZXad7JVMBBs+E79WINBWqZNYyfeOVmJqsJ0mbv3K9zTzGf40HVDm
uoDkPwSCMiDYpJhT7YiclUzCV80DPAod1ZyRiuBtPzpyG56MjSBysP9nXazgXrlEf60XN8QbAyYP
85wvGLi2iVaOHXBomw2cZxgdf7jkwtV83152DEsKVl4pq+kZ1Sx4o48WmmOKOty6Ggb6WewugV1Q
nmxq+exkkVckTAysmgyks8QIUo9vEl3/Xpk70MZD6IQKF6BbPa2ctqkzhWhyjky4Bx/X15ZM/HHl
BghxjGJTAOa4vPhJDmbTdBU+qMYpJrxtkZgDATYAG+t64zAPS/yn7NiKbIlzhfIysr5MY72tYDky
WU/SJv7b0j3M7CYifORh9/vON/mr0qAUFjiUTEckCVppwVsHtJ4sqtoZ7JXWzSmAbIDKfCUsudXV
5AM0HI7gaHYhj0xVVQbJIdWfqEfK1bCkhmzKybEK0l0t2H8o1YKLXonYdpvtoatfmR7V3F3SwKzX
Loq1k47BO2ZwWGkRsn5/iTxGBSNA0Gq1MMMY285pbQ83q/DIdEArnSxkPIGF2lLV9UBLz6dm8UN+
aR+BNH8Vy3hS8lWt2e4RRk6RI6TRO6HJgYfRjCw6M+Dwr0YuVzIzWQ3yfiI3D3owZzgmiroV9t/b
TXXzLq6B5RxbpqXdbZFRGF0B2iVsErFe2J9bbNGOqQnw5y2H00KoiYZkTWIi0nLmd9Mf+xRoLVdU
pJ+rU016uspdt4I/WOu5YN1tPS3W5gNSAcOzle5fbgRIx/TRz8snh632xbC2TSBFiJYJvSroiirG
aVj0B9ySZi1m9kIUeP3LTcytdsPpdIPRblT2x8QdRtpC62AkNRK3bpYfJsbcM+YBFXTXNpZNsQqz
priMZ52Gg0RO84x1+8WFNMANzuq/LrUkefzl692qnnuVipZjaMyTPpgD6FoaryunB2CIS7qyCn4z
xwJqbOhpiOoAWVXOaoTP2kROgcvlVHPvvqAM/UI5MXD2zsUEh0c9alysEy2zv4kBo0Bm+np+Ur7e
BWYQ4vVS0aIMIfEdb8cL4jsnh+yUI/zTOvVbaRj0JEvbd2+Qhmrv0aJlT+7ZueW4VphmMlcMSZXu
jQVa+Y+sHKisTK/G52C6jR5QOCPjU3MBVPnrvSxTmbe1uDj8r4lYFvBrKS/gOSMjwNNdRag/C9Y2
MAvAPbyRicfjvjovKhUi563N3wVj+YsToEs/ZTxV6Fbn8vphEqC12jf64v3hv/9hkaQ2S9LWa2bf
NYGxrXBGHcCXtb7zKVISa/H7zx/rduy4hYUXLxE5XTnfGaaD+SG5yUJ4uGZkXBTWulIPoiBK9WAt
rvHAASOZWhM+Lr2ZzGlCLxRdjOjlkjLxGHc5AF0mhJJKHstM3J9kfKhK9V3ObFhHMWFREfQmCpwP
AWVE1hYrCwQIB8QfnH/WBJ8TCjLmZ933YiF74o1r1gdX6UOnfW23QAdHdMpMsU2renIrG29jR1/7
nSHCmI7LImnugNlbnUbNuTQkSFV6Q6vROHATzTn4Bt0++FnDfMlznGI2AX7WOctxDK6aYqOOrBOB
OrTsOgHBVFkw3zkBhJd5SEZgurQt8eRV8rk7IxhUTzavlwDFtZbl3tq43Q35zeVRzJCVZ5zqogxB
mAJ9gXBgUXi5AhqUlQcGEJjwxDYWU4VIpez26g2MbcZIpoZTBhanIa9r78ki4+ud+Dw5dmA3d+K5
nHExhLj2Uw8vtRGyv4g4BaZam+T+h2jpeorBDDrZ1Po8gqkMYmW/IFjSOOS33zQ9yAj84Lo/i50/
yISWXmFYYxREQiKZSb6ztnijHt9Y1HJe2R0a0qrz3W2ZNvX9rPL716u+cvOc4vhL/E7sdRk8jfk+
74sVEMPYn6SSVcXj9zhEKdyBSFvyAhwLAVNYJZvm/mvqTME2iQ+SrITUfAWDVfwm3/xl0w0iQMLr
oRUeNfsj3SfYLQcRKd0I/trs9R8iDFHcoa7YCtE0QXAsieIpoGEozphbRWqrBcfTw5/GrNWSwwoP
/B9gKAjqTIlGI3ICVpDtiH7+ik/NSIoKHoKXZpWb9bsXRknlwdeS2paLkC0HMy7p1NzsfPfJllmT
HAQSTrPXtGCZSTdfAO099kwEu69Isi51c5KQfKOWPe2GBxDW2wEEpz3ARgFPhS1fHDYW8ouFEZpZ
MO9Iq+AriIwnvJ60k0htGznRMYgbCDQ/H5FXKSB+Gv3zBGhbvL5SmUakGnOnxoU5NaU4JDnPIkEU
eHnWTWrwPmplW/fqyGFR+Fc7voIt/GjNMybKxfZ9QlAMZfPqe6cCjHpFXXbGyimrj0llcsA7TilL
xv64Fp9NTihB3uSKyGaTLY8yB27jKspbiOkavrz98y1w191KRCpEFmFpuIs2bSBl+usqH7nld1Zu
rmMboT4H/P2dJ/Kluytkih3DqBPqjtBbqNtN18NxV3Mdo+g393OIR2eqz7o9+42tEWd1aF1coLUj
9XheE5I51BWtgsWYu0cxOuH1yEFGi6/nJLxgxxDwmOKpcQXhD23z36Tg90a0wp3Jt1OvZAAvjv1P
fmV50AYw1+JCAVwzh+qIyQ1UwJ2dzxAm5m5EWk/vAaZaJRX4fHv0+YnGrJJgqewKWbaZzGbhI/Bb
zNbmnE1U1DK9bIVA61jx7vV0tmfpKWVNSTOanX8KBhxMh9RFfUxB700VVx7s3Y70AWMctL6jfKYf
eYnQUAiT+O25N+xBUTGZyEeN2heP94M5I7C41lfKWssaBTs+v+Ia+gc9/Sn7lervwBWjSeZXPxuw
9e4s4bZaQkESRA80KTUBvIjTFSQMUBR+vY1oAHfZe74curtwX5ctplOgKn2L7CKGBuBnifnKxh56
65+l7ncVqAewrCfXaHe9Xa0g1OkRwg6a/B3ywKamAM9TThkUx1Si1IBFl1I+3rl5wWmz/PBXdkxK
E2XcsPT+OThD7xFhpV3gL/DFLMUdXWO3lr0oewPoxHWUsHNIV8gF4+1B4o8bwPS2z8HzCQOqphX0
tvsmXjtbd1zhd8rnaJf6xwuqa0ZPGDP1eqFoJpQ5FNvw1/FoUw1aMvxojZ0gOdxz3GNPDMzcZb+v
7XEC235vCEkGgunPay/WS65cba7iS+JCaQyvcRKijIkJUaaOqsYlQRYeq6su7Dso7iP/iOjVNI7K
WSolYB+HSAV3Lmlp2wAmJ6H+f6Pzz/vSMwdx4kazL/Fp8TwQl5nIB15TF1eZYnhsosSnM0Lp3jqm
/IzyqxUiCUZekBpcVDRC22J8rEW1LBKRbmZkH5ijjX1HIoYCe9TFyqvpAC0ShcE9Cr6i3OZBK/V9
PmyZhmw/jX9HZpDs1oAfWe9FwPhaFC6Ba6Ry6g+cnn+w0IzTCS3NTJ/3gliIjkFwDp5hTUFePIwi
ijWCgSJfrRdw7vbT8wy+/fcu9J90Z3QFl2xqaWgPfI7R7CskdUWwsM2Elvqwj7rRLJQQXLIJaszs
2pewhOHUPkyB4soWaGHIXPAbRBmKzOFQQ7sM5sXQgWxCWnF8uKGJ2HqNT6QlsmWB3YbqFPo+xyH3
jb6FFZdu6Eyz3sN4whW/46Gg/4n+CJyWxX/n0ovg6/Jjn5/x+Qna08Y+aakuTe90ARXwV5XUXX/Z
nKNoEsLN93IKPQIMbf4/KdGH4wD6RCaCr+Y6QZ0QYbCBGT3LzA44mtaYUCb8SncInliiMjKynKXl
ftXmsonkbpNc1pgQx45dqMJXwdt9qk2AzTJhGw5AlQUEq5SZUQh6VkukJVc/cC6pI+S0B01w1ouS
WX46VY2Q5FcDH28XDiDLbGhXE0hjNlq4qdiJD9KdvMmaPRIljLD9wiUhgnp/H4mzQis6vtOcD7rv
CXDoAX2ADkxJqHqX5QoCR5QXF3yxLBb/MKy8C/T2dM1S/Pmbu0rxBip/PU2EOPVYuCmB6NKQAB8J
+n/nsI2FJdTg7ccVrWWU2tPbyqG/zchu6bVh5PfYcUYPfbnMqvOuZJrsIJO5ZvmXpqgxVCtOB6fJ
Vhvpehgz8gv2nwaNnhm+akVKTw+1bqjsfdq5EqOyTxNv8ulKYxlUvQp+CHqhat83byLjpOBzsjop
7P4A/uUJtH9XmZGwwI7cYzlBleQsocAwwF5LQOcHWOmT9V/ur+0VQZGcolMV5JyjbNXd1ywLogUf
nz8Uikj2SLaKykNnFRyuOm1jT5k5sVFl0aMlvgpJVc4gM2g3aSZW5G0w32XDs3Xl9jexNOFLB9LH
VL18A2H4jjWXax9rm1vzn2ncVfR7ropmoqI6j25Ch7RVDQ+cHklvqEVPkhZeCMl82PwdTDTAqjme
LnaMXq4tbBle3/4C7JqqzN7ehAyRg8Mo8e4ThkAFp4ymDiLEn9SMDchvS9nuILyQH6VntBgLP815
hDW4nXijYNXPWaqG3xL53OUOL8jVHUTLKIfBqPXvMHns67xRtykrZB/pUSlU9pru/utyQ8Ejw6vZ
ZMFmirU/5RzCCWyQtLGtiqU7TDGOiR7V45PkFZTeC9mV5uf8s7nnGtq8SWb/0ZtUSRZpvzzzqNbp
5OUtXfMasEzvnJa6D85z/PQFCB9vjxhdP0J/3I74V0YxOArBM/RvQwVSgT01yYkWd8eEFX/nBCRs
x2c7rxrjSDgvzhkGDAwGhfEx0yXNdxE9JT4GpuldZihDH7UCtws/cLbGuROd6bIB6E3fVZPeLDmt
OxmYTHC02SzXg6q2it22yb0+o5aPmkHUzPPoOQxVAheiKd9cpdN83WhVGxwLCsKAdzwxVTbKDEFn
mRKLxa+RyjH01Q8x5rpFWSYkP/I0dflEyXhtXjeN7UtHncSOKxDuRwlkGLQtmMm1XZ7NeKyOmC1+
YpAx1o+I1BIms1S/uqqRJPNJIQ33mJ78fXCsEUB8TpC1Smo06bvOmZRULXzkYlyEVrZs0KNLH/Pq
kwDKruJMWkK25k3NYYNnZf/Ijgz6KxduFjSgE6Hnvj8tO9QK3eWaAsCoC182RDeaER8GcEWKbsUd
NDkzCgWEgsB0KZTo/YuTVzaZp+zgFSHYGifFo3t+M76953FeGkiWOw6GHBKNgKLOTCUOCgxJdbjz
QRGYm2bO9ymyLEqiMqXqoi0wuHx+gKVbdmky1u04ug4ZwfJ7cuY+ejmv9TWvV2OUOcT+rXEHKFcQ
6yVGRDBt+G0wI0boN0O5ictv6vEPTPyK8SF0i/FRETondp6k8adGoqUlyDSmAd2sO0Y3sGNF/PnE
pAEMddO5fi9mLM8N+i2Rwut+G+rmwWleK9jK32KsoBI45zxxa39yTlOYV7qZnaXo3AwsrglETTS2
lSSPMGeUHOBcuPRyEER35F1TonBZoDC4mr2sB/6R3S6AdTUnDiAIhNQTu2cvTqvl3XTdTTznzh5W
DEfnevdiOJ1gikRMB8ACLU/ejDZE67h+KS1MDkQrucxYgYm7ho8b2/OmyQFVKP720hcYde60UL15
ZR4QpmQ7ShtXZftiL1SXTbX1qCtRBZz6DJdN9VUV31WfpO3VZqsxquLu9oap8HVKTUiDkFdLb/5H
846whFy31u0Qz+MvKuds1IAc1RYO0oTtJBUeDwM081OxGKO9mclKK0XsCKxQPD14AIG3OKK4WDbb
9YBiPzRDOHcrmoR2iB9CFWpVBXyHkN21c5lYr6K/Z5M7LnkuU58H9dJJz5fcWgDYj+L0QZDqK5Bl
v0/SinYiQp82PXYSnqeKW9ZVZWCMPFsP2nOTU/uYZvUfXOaxN0GtWOueqCqGZ6FMmR9eL6Nccjs7
L77DLY89Xs/4mo4Mmh5TOHtfetHZqu4tx4KW8xzrY7bZqtti9ugAmWKfRimfnxWWDHyK2u7rog0t
+qi3XriCIgyjpeJ1lZ0kQeLdUdbdt11CKMKsd+cOGolkFrQGv6a7RAIlu10/CaU8HHShPwx1wJ6M
c79ydNsXjtpuIm0KNrGwpHeNz8htTVGehcNofIB9DRhxnOOZ99+kgIBPnCEEHg7bpYQbR0j8T2+1
+UNJpVEfx8n3DZErgjmbr0JB60nVh297iltel3vtPle/FZtpEwg8YZfccRKLwAS49GbyUL/PMiVK
oa4p05tUrZ1MAHLaEzCMLhSIQStDyduv8XkCtbrGBGJo1PaHIdoTlZ8wgou4+jCJOZIoAKuN4dWv
NZTKXshQkhutvf5tb/zzIpRo8ZI6OWoAQPNt5RP1wmk3ZmmHA684IPpMqNUhI1Tt8w+2WCSlPbTz
5gEKcKkcaR4iyRREOIx+8wD2rdyuSGP/RJSM9XxhuLeita7KPLrJZX6XbPS84/kPSTFcbnD146N6
iYF7arAuCAT+vlCso7Ssx5UbckcT0MtyAB27s68/p+Ak60uGsd3huugLvYv1OAwLoh+1aKTPCqil
PTKuBgTQplhU6ppkYPKUYtEE2uQvy+ntxE2BrQoWpGoXvwHKSuGDQ0tBTflWABMTwi1wzPU5sZwz
zZKXdCK1YC5vedzu6mzCzkW6zzxfvzJtKrbhQ7XpzZK9GQYqcHvea/798r0PYeH5RsN9nG7WZHwu
bwf0tjqAJUEP2EY2bE8xnOl6QaTbaRVjGo5nD0MXXvCTdh/c6SJ0C0hhOQqMQWZXhR+OQd7SYQv7
YKLZ/7r9SdOtkIMcnq+dVbwfvbPBcQe4kjpWmxKKwjo9I+c4As8Ycpkk51JxP+sMD0Du1jNd0wGA
V4TaaiIFQSkhRLaEg33lW/nhTeSo9Xkdz8c7db+D7NSBFFDqXjsFnUgnRXoNnHdvQQnu836mptrI
tq1x+u8PzY+rioqYLVqv1BvpevGpRVIURgYnkn+tsAzoDF+VsJT9ihTIEJJ8R3JqAxor4BTUXsig
f0fdjI/qgoQmcTbPP47GKiAgBQuVDekN2nxfha3zMuiW7+WySacMq/XneS0H9ZnHAtb+/Q3LJoCd
o1r7c/UKVC63uTsu7+eo1cb1UeZUzlR8/zSSynA6xkYsrv10ZvvCtM/9+MquNKcEP0SZfHGfk+Vx
rQKQTykvduL4+eUsbjJEJjeWf6SNgwEc37Y9yW0rXjjJK2HqMh6zzUSO5KMbQBe5jyiezsYtfjj/
DmSN34K6AZb76x/06Ygij/78QoQBqqAca2JAIClXBTrC2Fpi23W8o8F0u7tB/qGVU+Akam1zqVSl
pFa5lCvmvoNhrYCbEPVhcy1vViVzDMkuzhx4+r9xMnEYeQxz4bqAUK+vwkJ7x+UyOxGBxUaswQTr
o0/wLg+hg6JDB6gXJPr/TYsV908GmoNJXOfQowl2C7UJIPdeJAwZixBxOQKWDUZ+wipK2B1hMn7j
AKx3clsxh7JY8oqGNBxYv7P1W0FMzk+eZnSSgeydryv1r2VhO6K53RYSxycrlQjq6Kk4LNOLfVYb
3m1+BdUpC+h7fIs7FyjPiP9Yow5+PWhZ5+G81tBWJf5uUOECnI9dDQIYr2MIKaZlEumJTrmiy0qv
ZsN9/y9/EZJ+/VvHq96e7nPbrUTDzvkGE5Rr+rnY1RFBnEgnLscMABjMHUTipiChsWqzecRmY8tN
E0gyWnGliKYinDdVmnVKHAsRW8QIavKbL30aZoiePVy9oj0/OKLCVRrIFv5DYpbt8h0G4TDSMImU
Rp1ZLPGtviSAfNbxoJY/KaM1CJk3rMsOZ/dW6puWh73ph2obDbULgNInd/W2R6D2ePAFwQMnARZz
EzaX08TzSR8LJekxyO9jQb1M9mSyIhhzp6ZpqXqOgYOgM0IYs1Z7K9zdLIOKAD7ryKYudDMY1Tit
G++8Rgg4etHLe/QUuA+wHRt+aXsho9kimHq9zs/fpTgrgu+KQcUgKekU6/MzrsnYoO93SkrMZC7/
cHmEoAt0UZFw7zrv9Sn9AN3fKjoZ5NSmU1vcRdSuHE4GdGglSSLK1XrWs/pnoF8y8Qbb84KgO29k
Wj5E01wNP8RsfowYDR0KC7noGVkz2n08+/yfWZB5plZdaju7OBxObnYqSvgFhBhLJJ56vooP3fhe
98KplEAjw0bMijQpL3N/ZWZDbFxQdlVDyeRkz2U7kBzDPG7MadF4Gpm6ekeMt5JNWy84cx8JWDzv
HpHYlGmQtxsrTsKw9O1lprMyLB3Qdwe7cXNlEeSWjachfH9nz+o8OQWjCdWVDWwQZeQSIGw3xFqy
0zLzYMQqekA+9elsYPkjX8ZQCC/e7NAbhfSc9dhRae10UU3pzLtQPiszRDcaOneaQcXuAg/HdNiP
0Bsz8EwTGYDeVGkzfdID8Pd0lm5ZrXM6J4kZLgGAYLX8C9925cebj8IpT+mDvJcK1UxmKvtzBw8P
oHt6it2OC9N7lWK8j5XY1pC9pj6CKrCRvQzAeanBTYdNTQKIujN6cloorr7n7KAHp9pNOfC608/K
YuWpbxIt5Js0V1BH7w9PNUR87g7T01nOeZSJb0zxJt6FuuBPlS7cOxrylbZ3bqWTApyyLNoS9a74
Pw6MthIbQqNHdftF/UR4MPrPKKadsm+goJCYc6nljF9jfRddl3gcAUKHAud3lbIktsw7qGRwf7DQ
FRm6Z4c1bfM9X2WhvjdZpz5iZ8+FYHU81anYJuz9rKxWHNZ8vf5lcLkrUvK++p+qzaekCrqIiHI9
ckUvisoDUZeWIf7h9S6MVzr60OADd18zfZxiLWnV8z5U0Hp25X2kqlVyK7quRbC91OxIjLwz5IDW
V9rrXQ0tNDKNoL2PEgb9+pBqy2y9nmB+7FJzGK6ZJptwfhDkoH1QIohwStGYVC7qiH8qouf2fvMm
7PtrqmZ1yWS2b+tkZu0BZLceBtGVY6TxCztEituVWPjfHbbsKgy6YX3zp4G+sENmpLk9LPx/XaTf
mNpN/V4G+UpOVclQMA5rdYsL6RqBOpK1yEdWMvEu2p/cyauPGqn08OgxNOYrHlxKgmuY6w/FgtVn
RBN+T3HaJ+/V857QnhDhVoV+0n+iQy77kEWhW/hAnGuZjkm57JmlDYgAJvi8QgDq4yI64CdW4xZJ
NbMeEU2PbS9R8CTvYMgPOoqryDbE/qZIwTUnJQkPLyxIBZdVr4E/7qNf+DcmQq3MwabaK/FDKqmx
q1eZ+OtIWgzY24vmbwVm12VU1avFCORszrD6tjQ5JLpU8Z22KuWzlcfzsI8xABdnFtZK5iRihMXs
ypw6vuzgfFiUH0QQPvBY/q04NMvcGJb+HZLqeuL6GXbGR10zUGI1iTLeS9umLPvhlheIcUZBF6l6
xmXADaZWGJBQHL+umasuFtgMX951nkyCOP8mrmjzknEg0zsdoImshdpRuAGlqjYq7hEZvq0CH59h
BQSrBKGajD+oKQabx7tGPfNnicg4a6RJTTnTcpS4tko3KGV0Wec5DydTFrHR1lZviLRLO7uYVQqo
01GH9I0elB6/VWeQHoBmtS5cTWO8fuFtFdSSM4KTbZlvQbbd9ShTgPwFDGUuYyMHhDg7r25l+gKv
m3+kI0bhzgZofM5hvI40pYMf8Ntbk0ldyscFHIbZmPoJh6N91N3eVBe2bEaq3uvLGJVH2JOqRxfH
LqZ01Icf0kko/Z8LePLMEX8BhGyrEpJcOcXB66Xvv0Nlrt3yiZRC+obXx8yniLVkLmAP68NTi80m
0kiwAgR8c/EbDzZqukggvSVocOEdN1uakKZ+h42sjaUUiT8dksk9ixQ8C0lQHNZWodKKpUGNclT3
xd6y8JsUhF1YEg0FdVU4SbesE/LNvkM1g1Fgutf3pzBqG0yeEd+Vb1YcYyrTvQTcWqw69TzHnVYo
xneFrdRtMgWRcdHVmuKCT04YJ5KlWuU4fSZBgm47o5GzIGRpPgrPX4V2p1oqyBwpwF62lLp9UtZO
KoIX4BDuLCqTCKmn01HKOwR3KolbWShbQ2KPf8wCXqD802zM46WP7QgJjohc+/yya7SWCeHh64kP
oYDtHGH2GTzI55Bfqvfo0QSAy8bmJZohPhDV3eFNHa461RtkcvaPLdwiXxb3ZYk2PCF+hKilfqVf
Me2bjxopGSMc85N4H7UZWTM7wFUxXHyCVSp+g1YkuBkiMd1cDkizxkTQuPLLsbYDolpis+ffK6bq
Sw1ri1/NbzBiPq0jpMUWBzPf5YbMvwTd1dEodZBAzgo1x+JqoPAMX8wDl+Kpchx6MR1TKt4YquRa
ZIdZhdi8YrT/iiK8oROnbF0oYljsLvHwdk77bF5bzrUARjFTcfGH+kpMADXkyT/6J2kB8Dju+N7i
U0arlTtRsRafZeFJeS4qQUhNFMgz3RrO1wE48uZHuosw99GXZXJ4Xr30wa9+hSDtnN7tNP+WEWaA
FIJtF2vshPktGbB1A3rfw+AWh70C0zvAHW3ZcyTWmmzE3cyCb7KIB0j39bYyt+8vGdLa8R+/s/sq
7LfLus0osDEWmFHuN5CZayCTx1ixy+isZ16POErTj89DhfZ+TGx5rsWrLsHjuH21jUj/tufr8I/C
oQCu6X0McssOEt53S/LjlxjbHi1vq5+oTWgPp5pNCrA5BgdlixmD7kl78Oj1RDz6kXQ5654hMI1c
sUrBZwfcYx/SCkUGtQMoJUYV/WI24WiWJqFoUV9EerohuKQzj0zebalW91r9MsBZ7RrxZJPHBBM+
TIJwc66F5gN0rlvK2j8+XmG69qoEYFjvvvU3Kb+gKYiuwqyo1n+XT+aiYzlI8wNwHVsZOAVraLWV
ZDtu4hh4IQq/8lAf2aX4n6krCW7fA3FOHMiUsxcdGKZIn+OA5QW4tBf5AkDXaszcHmG3kPpkPytB
2j1REyd0003KOp5za9OIv7YYSshwIgNMhwL/1kuEqnavDS/w0fQxlSgL/RS4IimXgKViffoWHThN
1PICWFATRT6fsQ3doVvmfw6my3YsYruoL77nuo7fNLqvNYMtKMcrG70J70Fr9IE+Hr63yfTxmdYc
0n90nmWmy5h0MBRFSey1YrazLCc/cteBAel1Hf1SnEBFDUeJMvCIxwzIU3Bf0V8BPzhUz71hhJ6e
Gi4Gp7hdB1xQefxDU9qEYLLESYM31pJgz1BTi/mQP88dQRjI7aNrvtVJf0Q37rAPZMPeoFL0yRUB
AcztjbxHLGTjomsiBFETij1TNujCIsOgvm87G9UXK/9WTlC3Culzuqig1Wy4zXOs3EG9qtaNxvW7
6o2mTY+RQk01tllataL1Afx4CscLq+w4by+7RTeEyW4J07O1n9wthODPmpRzPbJbbvecE4qZ0kF1
3/bFAv0/CEnLr+IQyaV2qxy9QhCfOAEBVSJ/uGVlWktAaQTfZyj3AhyIIYiPIN14JXth7WnHIJqK
LD7dFJ4PnbIY1heTngNVDxQ65WmYMWNSLWBcXshok/I+8BDuthF0yR92jVCLk4PxwWQJugEAOK6C
Qunc0nv3Al13pbU6YbTue7RvpskRstgco7cWfK9xtimz2yhcpvhOEKQkpp2bobaYVCZnKfn6EHfy
Fkb2ehhI4aFB/AKQR2Y2y2wsTKpq7vhtYWSdgAIvXmho1rUW0kdN186IPFJunIGtvmhkiqOdTSqp
qLVntuysRoYhVGjC09xbPKkaL+jAMisk0M+Lnoz8OjIxf0FiR2BDa1n93UNv/2A2y7yuOB1pTetL
M6u6bgtzCFQ3BBYRjWnltG6hfhBUNVUavwR7q/Mx9rFpkIOKezMFCqmy/C+RofqK+/chgE3zppP2
Oto7OzJNBKzeGyLebcfUI6MgXFOyCGXD6V4/1ThicmSkOIHs1F4umyUdlho9bakcX5+VQAjznb7y
avIRqMPbNR0zEhY19iXcN0z2G6FCQ5HSvsfvIn1Ue3B6YqSc72P/aszGtQ4Nwnt36ZY4x2yvyMrO
GfZWO54g+R49pxm3mCIbrMpqqwjUx5UdQtQsSqwBWyvTBA+YWZJ4D1grblsxbmexjkZp8vZo9ma6
OIv4z20U8htrUJAOAudwKox1NtlinrpZcEK7L/uLobGh4OvHHd7jfxxxhQ5XI5a5EAjLzE9iZAw0
LQqJpdYXwO5b08WhTtnJg0N4aHUpOUsPsLCKegAkT8wukdfZ7C/+a51CoFmOz32/hEdSQIszFL1p
7hDksx9nLgY+BBW7piRFx8pM91Sr1FzTzAM06XrjYHA1skx155Pqbl/aYLEgZpZ+aFvJDPY5Vowf
BvcwFSupV4MDY5T2Sa7hs83uvitEQ1fcS6KhWnVgpYhYge739qVPM1KuPrKLryqvUoM9b4FswjWs
O4AAGoTvxQ4vARodktcImMZhb0poAYG8q4WWzH7B5lQWnYRFSQxVjOzgPgWzgm2/AnTCRsj8LkGO
BYh3nAnV5t2fCr/a/JqOKiUGs7ZtsK8olNe/rpHLlsNFlqXIXVbrrtDTxK/FdUnd5hSO0iDctq8a
IK99lQwmfH61wc7mDS00v6maeNccPN9yfOSrZrVe+hvEBL92EiDPW+7MqED7QWBdQzCiDw2ldsKn
mldLcB8e6TqRlobYTr3bKL+KYPXjj6RXCIKK4cqouL/mdR34aLa5ScpQt+vvikEGIrybW0rtmbIH
fIxLK6p4TmCha0cS3PM0NNzxoO2RoWFpkmdN2PjZSOHPn1kVGoqBz3dOv1yJhqRecVB4P/ysaqfb
/+2k5RKwpK/WY1CtysYNCPwh45NHg5wXCHlxocbHuJ0paZtMfP+gjQZYj+1mLaz1ltpF2n6myace
0Cbd1xjn9h73+ZRvv5XpQ1HbEe+Kf1bhnlO+WUg5XPDEwwPonHMmRUlx261ry1TPCNGAZNl+mz8l
+0R1LdaKC+tZB0qwUX5+wEEbLG4vJXueQSqOLYXmQHTi6fri9br6TXew0NIsUfcRU43FJW3xEc9x
xdTX+Fwyz/JXoPmybRZKAvOG53M8xlfJ+v64FN8qzzidqNx4ZqahvWbP4jLFEypTiqH2g7m4PSCR
jeA7OJp+LuMye3OzrSiPgRF8+twBkZfCOfrNBHwHtMmJet40h9kkDREOr8XnlJOHHdjEXSe9ck2O
PXV+eUQBUAB4PhLEDI+tQonuxTPYZ0+0E4q3SmAcSJWakK9PTKtjojuQLjWEmQKCoCzb4Bse9YLL
Vd2BvKzpOWdnOKYfswOGC0B8izFhXCxWc34QI7/4LVlQkwbAcCXNtDsA2BdIF8Uw73rEIUxhzsGA
nJKB6KvZfXsTKdxcL181ML+0qWhBjTJFhgG22NpeqCpSR8/KJuOXboGh4fIb3os91RGwNYrCn2/o
6OEgdj/WnXcnbEKWvELY3xmdvcBb+esH7ISbHbZghyDwd99mXC0Jiuv3k2no2XHn9MeH3u9Ca7FN
he2ssAm2JXOAW9jzv1ksjK5pCMB0dluvRyn8HxRfg73ciKKN0DhBEIVwn/fEri85uDpZRNY5GID3
wGEc3ZhSi5RCn3e3bdbumD5hxl2wv4sbn+sSAZFqfwB326X9M20K4QwZN6pjqYqF+47uhbZvWUOU
afsrRLn2jYdvaubPE2O8uKP/+MGW8lm+6DFveCK7yxvQyGMc7ySZoE/Kt24I2DYUxO2tgYZvBK/d
IFImaEj9n/ypzbXqID6FiKM+MMb0ZuOpDCQrpspf4FVU8XG+CN+LF65lSG/VzG7pLwtJLJO3JRaQ
+IGdo8BgHcUpSr8f2ne0tmJiy6DrX7xkywmI5aTXOM6CF1EKjWs3a/9ZFfZfhjZruJRrz8ezfMp+
LphpNxHOrR6QrPZoYEPUeZ3tfbfp0K0GZsO6Em2+G3FLkIX8OCxhghy6em5mX6JiMVCz34YmyuS+
RT4ZsJRaqLTZTlQXvDTHPY1t1BaTKjrk0RBJgr5+sxmEnZ+tXgOLDFUaDaaJMmzAFNK2iecmnt/B
hUQWDp0blJnnuGbQ4dVxsPXUAUBlAhLYR1iCYi4XVNhXfzsVuHpknpwcSPyWdv3ownzTLDKaZM5C
dsErT6v7enxxzS7powj+T/T6+EvZgWwW4hWhirWvxBSyNGhsmW8xvfl/LjvYwqUXEGL1uvZXuhrq
8SBWpmV5eYJkwey1cUcQRq1ptP2FsJHMDn1SGb1aADscq5l/8ecK28x3Kiu1bDmO6qMpDJOfu/2r
rYmLPU1ajIcQwV99jL+KANuCpTKbW08hAQDpVbue1BXCz+y+nCoYYm3eE+bCXp5ttJqN8dXm81fJ
FOeJa8slLoBh5aQDsF9zMSua5N6vJsAig7sdK2/eGLesbRAPIiwacUMio0MYHlYBKlLzSXuRICTH
txkvDqtvAB/tX1WXCx3CYib5bS3BCuX8QaoEUZz6CBtCAauPUpi+0gAm55Tbj1zxuUz1yo3SmA8X
MspwUhPrY55ajLbXjYKbhBARagSbVqIROK0C3+GMDkGzgdSBf1gwtyp9+v23n3BgMguWJUSsWH9z
vWYrw2iwzM8wcmTf63/Ji19k7lI0JqVRjh/CbxyllPtq9w64nGTgBmF5FmtK7xM85N95qJw8aMzg
CeOiOHu+jrQPhT02G0qVmQGHHZo2vNmQDtfxTgqLzg1kYKCO81aSqKfjDe5z0x4HBXgg2DOH96AD
z5b9xUqPggt9TTRqKezQPUQRsfTtPvPZukGwXZ5ldGbGXr3eiGJDio3Jh6iy5dvCddU/YeGajlKU
9NaWinjrqbeIb+hK17ixE2bRnEIq9AAiIKC7nIocga5PndZCbI+ST48wjOmh7HsCGj9yMwUUIzzH
oaDq17dQOOvWPlCR6rHGrzQB4mLp6fVapznrFk/zqw7BoMqYj5J/iSDmQYRoymqk9xAyRSVQlub4
D4mgDA+8sZWQHsmwF47rSweI5jer8YxnjLcb9PcYs70NnyRqLIAoI9sgMIgWMXsbNtjMWJ4hT34Y
3foyhlzndk9iRg7c3M/0Dpm2JkjnQPk4VYzOTtu9mOK4/YRpz+RPA8+DmBbwT1trmPYkJW5cCSC/
Cff6dAJTn/Sdtjta/1o56hSg/suMVzp7vVXStyCQN2HRDY+TWqyCO4x6sqDpo1FXZ0+KWYqaENBt
r5VIFzQgvkuaY2z2l9SziZRVo9SBKAc9TUqOQRRZHwUCn4gOw+R8Du5Kk/3CfPZ9VbZVFzPqOOPR
2M0OObH7s0iABB9tSiO3TctTIbEwtOL9fZA26iSzvWhSC9zvm9RorGZZuKJDppVlwbh+s77QdGj1
ityLI72/gnqafXCIexlwFH9AmfShv7dCBSpK6LZxzY4NEEEFAtcqRmlEiLiaG5gL2tw/OKeectcv
SPVZBeVE9GCQpkwml7BfFoSOkXxj80IFAmyGg4TwhXZHJ2KCs52NuKoGQUw0GcPZsp0zi8jtjs8G
gXe3XePUSiatO/AF3shoaEzD3ngkR4zHIcbscayOm27qD0m0M9H6kYcke9HGrYtRQSkw/byAT6Pk
pEHvuWmOzwLlkzWCNmES9Z558sUoY80bQSF+upWofBpHEdNdMKMNrwVgio7njUSLv+71irnKeFEM
E8nPaTD8NgJC6pWBH/WhvvHLsnwC0RgFvIM6pP4JaKUyMYAdobKN2UMJT6/CNLHErGbPKa55DGX0
jAuQCx0xBMLX0augyMtipsG/knwVymFBXEpa2C3OdOB/pTwY6hjgpoQJA/Wet5cgdjK1DFqmQ+vp
CN2E27WldWrWyr4q513lTCU8tUUHTu3z0HAVQxzV6l1J2heiD/22N71qsecrdRjOyYI48eFxC9sS
DHA50j/szUFOMm4Etm8hm18B2JQi5GHdukZLF3LzWL2k0DJy2EAD1Wooeq3IbqberZo9IEsrsel6
ch0LoQ8thn1/R+F9bY6fHU+WVOrGW3vEZ5dacmjuK17tsNk1K1dRAiWr0HhFU1K062vUxNeVfo4Y
CLgoU9qUKIwUZlxZ+GC50xKjS4R/JGZVAcQ5nFXYIDqRNkyii43CrPsSMO8Lddy96Qk29XSW3z39
AAMY5PQ8WG+/hBLKBKXnp6+CmQcEpphV2kwy+k6wS5AjVaLH8CyZc19nEwGDKVissZU+60SeSHGB
iLicRo+taHQSx+v7Dzu9qlxLA55+uiEfkmbH6qX1xkJZgCP1uOH1PxRRcp3B+6Xm8u4iQ+meo/Ro
c4dDp2LgOZBQUxZ055UVNZa8OHjY0jXvpIuK+OYSDnSab+G5vYK5lKPZZN8SoBIVJabq7LyIRwWX
vbpmUWh79POt7AEUNbHK7ralXJSBy4XSrZlsfoMFyXJGqyimcJYbZeHP1QyrkcrPhfKHK6lw9Ige
7UF7NTejK6esE38fuHWubhEgb5dtLNUxjx3jfqbtW6n/ABt5s53+p0d2vemVkpa5gHHgTLWA3FRH
Jz3rHn0uJV1bJyiDp08z/llwWFGrXXgSkeFCOgbHHj/TdAvt+DLmskbOQxNzn/PGQ8cNvvfdPf+k
IY9iA/SsvOtL9NAp9NuomkxKEsMwXX8KIs9UusS5PdeI70f8t56HPOT9P0ylELq7ZJD5JCj/h+fK
FFRgSLby2ziiS3JRtIF7p4IbS+TJ98tFbbsz0BuKwBD1uV6R85N1p3/lO0dBwirTKzUsXqjTnNjw
37BauN+ZV80fCEx2aROmNdfAP25OAKOkZ5bA49kdmfoJb48NZ9nEjjsH/2FvrWnu708gIW/LG06s
PY8KwFmGBzn7VKyyF9Yg2yr038B7iouEU3huPUiyFjFtnOU8OrHsKT9HuK3qubJEpsqIt//52ORV
uvw9us/PfircMDnTnANsjmLw26a2KSpXSNCy7VgiiT7ERPpzi/qdulg/hfNABUHfpBTuLFZ+UDPI
EtGNF8WBR+vtUEMNLYBp2+GlAh3mIT7kupfMyqSIQAjTe1WAGTVMbzDBtOsw1NA58J59f/cW+7jN
ZCVgCekzbsyRLMwEZSepKtvBbyLut9lk7GMs1zU4b5VXZqtVWxbTsRAkSjAyamXpqgTh75nT7FKc
835NtEJBVjr5fj7e/jlz83Mzvmct8FdQ7sO7iSvwegdZSQwiiMZIWbRD1xvHkFM7aurgYoyLPyLG
LyBID+6NgrhqXgPP/HnfEuvDwfPC7ctQ6t7Zcun5kbq8mdvelWpHgNL5AY7LBzHVtX2UiB6l5v3y
ljrRJn/SaTegfZHYHZV1JCQwzK7veMU+miGUY4XPhIduECNmh8RkMVzADDUdV5hJJT5zdhFd4KUb
Ng+JREinhq8Qy8th/KWdTt1OE5N8t6S/oNK0XYEWFCpPqtXtZ+HhrwuwOoPf0u0hEIRILs50vzNN
17n5yShRx3NgplB0gG8sqMqOybu8GNCIwRbAJtl/lqkzaO1CvhwJfFQdz+byYCGrwe6qZru6CFM6
0wHtr0NkFEaadLTEJc7ypAUJsAypsdQwm0Al69Rruje/kYb6u6KFwx9f5f8Cq6FSh7qdaK4H4cMy
jFwplLOR9zVl5uRQQgW9QPQkNvEffE2Ax5sA0QdozbzmDZ5fp7yfoHsA+vRwGjqJljjIG6sqcIHi
oRpB3v9wVxe5Fo0FvR6ASYnEXgDZ65RaqUThG98Zbx73rpA3K4IunjngYyMv2X20qubN4QlepuiM
nVMdvjAGuhekaScEE8j6AWaaS02g93X60FwhxadmxCyD002eO4G21J7plgjBrIYl2BHkGO4FXznd
74UQcUMmmie/TYPOKnlzYTcQqRDBA98I7vGbqEVPgl56nyt93VhTbY7RcDFOILwJqOheif72j2i3
N+v5tX9y1VswpdP4wOE5KPPy1721cLzJXL+R1dnvrYsFlvCnDRg4MoeJ6Jk6m4+k31/lqSZCkjYK
joCYqqIa3rKlivkMmWo5kkmuPTjj68dkiI+J61/uSh7L+/eooLaQyg+Rd4bS7BDKVwKyw0geYLcl
eOcSqRGCYsy/02tfyeTomxpMEY8UMgB2s2KPEEqiTMHPVavv624QKFoLYqaJQDXClExph3FGRW47
ThYWDruU7DyeBcTke6qNlopwxqv3077wOX9QR/zT0vgrPiZPmLsmAwIZRbP/PFo8DDDyVdjtWixZ
Z0GVAT6SfaeUUmYuOn5pjQhDesA9powXItG2h9luxbo8RcMXbW+sWTD4TZsy2H7aMWvveX2jKskx
ozjxsrvwmagolmTkq+0pAf22l8NQzpqDAEmcgWNQ2DyfKhfNoiJRJmilQteUUiVbtmWqHcLYALjG
ukoWQfMp3vh2zgq5r+8ufFl5tVIgBvvWEa+WmDxrFZWAhOcCOnQHQ8VOuB8gmY99cYqnDWRxIn1L
NjsrVjql29taB5O3zISH339KHc/u8FK1ax37uUtPABjNdY0nGoc1mzbESWqIINYnvMIgLCrSvyqc
raPoio75DPPszFKjZe9ItFuSvVxNr/tLezRUviL/eemvKP8FApcfIVxlP7BT30frF3OlhgvL5C0u
nRTTMSnIXSwd967+qKG6Q6v5kZ6trhpswWtr3KmhaiAZlVW5su1amsKfX5QKSqRDRLQKp/JnDUjw
l6WnaH2H/Hnw4SMUenEQwm87PGiNVlY8XdcnviY5uvxs/oniEB8+lnrE0mUcapYlNE0KihV2b+Tk
Whnl609Iqb08rrraClAOE+yxVrETTF6lpguKmL7ptCPJeLcobJO0t8KcVa4YEtMMwBszYpj2V8XZ
iE6FkBdbuUi6nNqvRxWE8DN3tZFVqcE5g+gnksR7Z5pmKf1VjrzxNOnjHACwfyZRxpMrCu62+l+W
24rlFuN53cn7pd5hyK/hTt0LJhRXbLxmzZM0huXcFc8xRkF70drGmBKzab9Kxesd7oHf1t8iK1H4
2HIfjPYWACqmxdC5SmRUTFPEpskK5krx2QF/TI5ovMa8J6u8iu80Uo34IwZjeYqJgAsKVAScdhiZ
1dd9XuWuMNwRAFF0HxNMjQtc8RaOO2WqDHq6z+bkCovCi3pA3sSPq3jM8Rz2akfUD2F1vkaMYQQH
8vMYRT+6kU+lc+SzuNNTTV1AdYq35518ItnpIDqE98FnCnxG1j7vLb68HiYwwhBPAzLVHYDS1t48
ZN7pc8EWCXoUhzCOtKCWbwuB2+pZ8VqZ8P42HkrQxFfZE7BqzBfASOGGoeqYFBd+SJ2NO1FCzQUf
XIW6vo8R8VWhRg8XzOgXsRhb+zstiqDoJzzX3UpBM0W4zq45IhF5ojR6Cht5/w0vixmKkRTzEknh
HnH5+B/Mt0yRWSc05RQdSGjdPsYqELwZ6wWcW5lYgi3NRiBtR05xAKbTa2L8+7ReyQTC74o8BABW
CMZse+n3o/3+oGYMQpHZDm13Fqs8xtSJLMpdPPyyArlN6Oj0udQ/RgHO7fCKO84ysRcwZI95LQcf
iMUmI0VLK6zcaugGWAvwLaJKkTSU0jFj5r/i27oqJcUX1LlIHgmFIPd2rmc+Om4ZzIzFd7rr2ibl
a9wdaTkpxFnRoum2t++y4q8WUDyP5DTGeh5EOdZclOz1O5wRTdPPVTPD8Rtg9beeGHCumGSorYeE
5af8H3f6mbzDyzc+zkxj6J+sSGR8uwmVzDHzQ+zXEJ/3x2WK8OeGmP7u0/B31lZO9XCQB9NXUX5X
T8Fzra5sPnY/xxNQ5naZpvZNIZYxuWqXcAECE2gk+JhAKiOn6M8RjLHyb9VMU5GQ8XuiT84yXu/x
9XQ+GanNo1XSSt72SieFWnb8VJahtC4DeX8ysSHUL0RVI/+5oJ6EIgamDSufYy80UFuoMFVskank
R3GC1szw9011jAqp9WqtlFAAeL8imfWlnpnXS5EfRk5FY5Ib346KYBmgxf7qfysMFh51SjNjysBN
MTbHxZ08UWTycGdp10XXvXAJK0VydVOF7fNORIEpu0Zm5ex5LPEhlQBZrxdyp56sdjYVduVd8NAn
HHICb9X43Z/0HCGp0V7vQPcxe3Y38JuBCUoxWjQBJjXQNrjahis4fjD8swrwMSrLex4/VQe4FO8c
OvCLI7Ck9COdc8jycD2K4vc3wbaq0VBqrXnwDoO1JJpNPiLUuvLaHz90xP25dIcaAGv61ddCS4/3
NaFuOPN1OZqw3MUFqdD+nRm8uN5sFXKuJHuBuvI57KX8gHFp3WmQ84hvZhpEoAabhkuqg1lSxZv5
eNT3FIgMmHgR6gROxLahTZZ9CVBLMc+n3THLMCiIirYHUdNrzkPgLS+78SAXZvkh7CFr5sGehnBA
gAVXWHzpiKNcz/sLVbO7jhvjQbHIgDc8AYkReHjXQcegZMTbk+WExSVvZJCLMzoGDPCz7eAIdO8/
4vJIRMfJy/6roD8yJesfmQ+yGEnndMo/qP1NWw5E1Qkc0303RAJTsEhcFbxCLrHhp1QtGwqgSFJ+
XkX9Zb4IpJxf453tcLYak7EqbQjJDmIOAor+ZUBW4ziqkMz0h+Q2qUQiqwU94zYCmPrAxkl+CFdr
h6ECoILqjDmkQa0NHTWKjC7CIssfRUn1+fTU7zvh/A8ImbhvI08O07U3s1Iotrq66AN5+6rtvaJV
JENq9RwANwFtjjoOXd/N8AWfEkjkop6z77fRMH1bGb6UQUONVSbS9auETDEj88ZgsGfa/m4cQtiy
yyfXBNGAPVoscYBMejHxApcu0Sk7nFGRj+P7XEonwQ29NsfEGwwZm3Tri4NxRUHU6dEdvCDIj27A
Vw/R4OrixGmCcudmYZMYALIMaJiieerJEceJ5VjbfaK6EFiY45oooBQt9NANzLB/6PiaLlni38tv
rWaN0+MhrvKqsUHL+k4sidWoJkgYlzb8v3HqaMc6JVfxjD1h+Bhp5lif4bh0fZqaqYa2hsXlD4kC
g09LJDS1GC3jdrKJBhcFEqdBk5ZjaS0E9Y5BdzGfnZtsBBQNbQz7i2es2Op3zBJVeyAWN2ICaTEf
paM1g4+vdcmbn38kgqKbBnsxl7G5H/nbpXB8rcLVKAHn/b6sNWL/q0gV2huVT8awzbgdHDoVj7Ry
ZAFk65wIcT4MJYx+3hHsJoz1GhKL5gFkAM1sWoCmAh3jvpStMeq0nuS/XedZ5/AW33s234WdL9jl
ODZtLhcQOa4o7PPO0sSfZ+fR2GvHTor3uNE/AlnaOYeXQ8dZ4cJpk69zKTfFZuDX5Uq2o+WEWex/
nL4MoggAMnvzD8u97Gij6VAsJLOZdx39i+CYz58vTlvvaI9ZeTsF0hborI1kPcMmMhTRWiJt9XOD
MgyLMjLJPdUyf9Qcuqt98n1egCwM69R6KzY5kng1jE3rK8YEQf+ifX6cG73LQs7f8hgShnyaRxnI
yfXKetcOoUejNGKegd5GsghOy81DOL3SJksMuEXBuU9WW9T/DHPKg2Oa86qp/13GnzAya9bsLpus
fhESEyLf89TROjgnoCUXZgZx8TnhRPaVUEdGvGwea0U4ZhguyD+3T87F4kw7mTiM/iya4g9dM4ZE
iFRd+CL2Zl0BJavr/9Iysomt1FYwicaN7ySbkdG3qTYhwgoYeU9ARp0ZqUXvoWvVz5cYKCRWUNab
liPIMSwNd7hszU9BuwdBLLDrBnsp4C6T4lL01Feit71bwpxZ/gaNDYLh/kt6EflYXxlD1ssjCTur
5a3WBgBkus8lsa7ImrX9QlhlHn2UlYxb0j6YQwc6nz4JsyC1oDAqxJHGqU/SUBx7nfW15XV4PXUS
hArnhyBPJpuEsl4CEA26gJhu1OoUQUGkFGwZkDIu2Mtb08LN2yylubd1P8EVEyJ7Y0Wu2iO2z41D
7H/Wkll3HzJWBBOfSnxLDcx0d4HSh8Xb2v3lkFPJpxvIvxCV4Qzc9DEisJ+3/W4JbAvzaYbC4I2o
FdupQTaVBCmUKD7TV20uqg33qS8qZaao833cfEA/nE/+QtuS0q7QBoJyrReGr6Br/ecbHwmuCQTk
M1buIv0dCg4yhujx9fARznKlf2jC/BYJOljW7GerSg7pCScIcsEl8hGktFpl6/XCdtm2hDHh1534
KUvoaVOYzJep2SMzTpOURPaDg0oQs3UQYcETKC6AOOsfmTGYc3t5dSruwqh/X58QUGtcIiY4WCFd
jbs+i/nI71KWoFLnTesCpmZYPcrWCy7rtNpnu2xDo8TMkR6iD05OGKR06QY5mPq8DSu/MhsJYM5q
lm3JhBRDYinnmhcM/VJH5gynrxC8DYb2t1CU+iaNJcTAsYgxOwscMvP8x9sLgVD87o8uWBAMTni4
YNRs8IVjTTNT9YWsFQuvG+7AKXc2lq5YFUaVXfRV7ZhGUZ4NV0fIQ66ac1gr7FdypDIJHPvlwUXY
2/V/QsrpzfhXGfesTW9OOlCtg42w3a9jXUtelowFv/5HsfmaVbUN+vSpu2a+aZoxJ1ES6MmIW/3/
i3y3THaJdFZiGQlwA5fa9bIkaaN9iJ9xNby7flY41zLg5eCTitrfaNvmxtujVmdg7uogvtagxqXS
4P3ed8d2opdPjqi9pSbs1csGm7xx8i6efD8uzbg459wW10+a1gX2GrHp5MutWYg9t2lyZgcYVP8U
NJ3y4Jyj5Lg/rHD4hEgLjYbfzykZIr7swq5DfrjPW/HUOvFZNEaPUc/wdWPMgaeWA2WIX7UamRKj
pKw0nGgOanTUzy5H4Z1koF5R1EkdVlGZu2mNzFeIcFMxuNwPDqSUJVM5Q5mhbdj1lp4aOzERQ/yM
qlmdDMT/KsAoIqVeauXiS6CvlF6h/O743dGzLP8HofAS4pSBwQO8EvoyFcqYjJSqqc8AmPuUVZfq
wHrQYpK697YNThGfspRTi+qdGpQaXxb9Y1EeFH2iiBsHBbTmdf+vvtzDV9fr2Jqouv0/w0Ck0VEh
fXVLxC6dGGAJlEPrAuDJFl/ti6teDufVanY0HopAcKLYuV91nOMULQGdV1YPXEc0L0vcT1PY1pUT
Og9mFaJ3YGXpRxmULP6KTxnZ1teuP5ppQbEyDBPGEPRvjHQSm2LTTC79pEwtUcOfKBI8i4SfpSun
NczRLQ44l1Yeds0dp7lG+6QRMqjbKVPz/0wE3+K3Ooegy1CtVJ55Qb1AM80AOOYsv7UdW/k2Eua1
8ADJdbdhhJY2mlKjy04HgDEJrq6EtlWF90AkcZKcpq3YrTJgiD2cYUHlBi9QUPUTJdrq1BTzlCYV
DcazrskWukLz6pFCHuoXGLR5o9PWrfl0MZypfLsXmO8aP1AXtv08SCj3TsFfqeXttDefqospQ2g6
CSkDj0llXvu+6CIuqIr8AZb5o9cSvs8Ja8C0CU8o1ybGVAFySOX1N8VZK6TiLL5FFnrm5zvwNWQB
MuNniosgXbeTZoNowow59Qy4IPCqZZ+AZX/e9z1FQPjpAxa7mgLXap11Q6bke6GgkFxMnq9xio45
3jdqU2BcdDJe63DxLZ8mg9ngAscIcP54ca+BJnNyq5EBWwv+rKRUdti6hs9aXDaIQbsWu/2Uhrl/
USmaR2G0fyzQBnmKh1yjCh95/O1i+FzDBYWE7JhWyKhkw4RnAmhYpK4NT1cQa0mCG8mOEwtOaGB2
M2QtBHwA0QLAlGfBksgC0/7411+GVbG/jgLqIdoz0bzpYiSKlmF9dxsX8f1BCNu/472MWYu+WIzC
hTwPE/B/x+/QUcFn83z77Nc0xqRqZyywOBC3ZryPzF7i5mifvm2kSHprWRk+Hodl2vWBBLUgT9NS
/ijik3/ffdCTdBanAHBn46tDwH/CHKfUPFiqQZbtvQsO6wNXSI99C75aSSPwyA6P6P8T+W17pAZK
T7Jl3QjSTLwLaH05kAJjvWt9+y9vFcekCDPW0dN4ec2+tJBTaLXE5RpKTnZtFGKVVx2piQ9+I8A9
NQmgjtNyefnH7dcIruMgID2VaiT9XIPvSkBoKTiVV+SZEE+dPNExMH4j0lvi7XMky71NKUP8CvIG
0pdxy8ipJcHj+IDSqGqvtVBd2J6u65toYL/h/G0iQlp9QlfSxEbVB2gORHOw58Opx3cuAxIh7PPG
vfw7DX0QHnEqyrbSqt14bLEQTp7jSi6LowAQkfTfD9+F/7SSDvCKT2XFv28/yxTyFmXROSQQdS2p
jphWPjN5IZYPfW9m9L86FytARG2IN96WX80vOuPh8TDLaimHIPu/p2PeLfqNJE3dDvA/Ihl011sP
la5VwquhsEyHbCAzu3a3gXYKpbWEgvR29BBinqAXOxcfj5i38xnN5st+/eAjpX9BMjcIL0Se/061
EpCBHPtvROp5B9xm2/CnCw4xv51DhFDnjorl9enJ6rGvono5+tunhZOZe5JUrdLltjAEr8xxOB2C
sBTIQQ5lEAeA9i23GDiivVAbhrL/DoithJg8vyykwYH3InrS9Y6UewfPxtcnajgLROBhnoXdTx6u
2xKzq2IZIbg3OO+YZRcyckdUURTcNF5LeUmILqbbB0EoUYtyLWFFcZqEDWShPQU7xcYVOXgMPryg
rkqJkvDi70E4g9Sr2ZaE9wkiuJGI3FFmrOQeDe1u7+nhXDWnfQc7Ye5/wviO+r92giMNdVj6sZ+m
yJMRsd6HcWF7dwUWWVGew0T0NdhlVrRhpr94PYt1d5aZzqa4ELRluq74MgUvuqFaG68rrnkapHLX
spleUrU1D5W9Enl9qJNYOlMEEFQY9Dxmmtl6NdIEWK/IX7o1ujEpm10i5MA5l/XbRKxQ28fNoL7L
OmbkJRjxCL3FcFr+m4OLLos0NlhaZAM/eptnp4J8Z8uaoHumKBf+FymUVS9tzH5zw9OMTtJn0EDl
K9460948dU47YrcUFS6jGGUqfv3E7ieDafRpsKaIq/BMgJ5wAUi9TB1UCT8TutPSWOtkZIGLlnWG
+CejBkGbTsOE1DjMiIa78o1N1EnqiirpET7emRnd4Ku6VmonBxWhBgp69OpybFCDFuuDvmaMowT1
MH8eUhBhwXhMdjG6098pYNnBsA+VadGIluBJa8Ry9CKTDVr1mNBHufUIi2nRHGPPF3p4gRmINiP2
N8F5KjtR1rMd2u7A9VXN0BGYdQ3RPg56ukl+57ksKuWRVRseB1sjfZLIMHk8EK5OvjCJRYsv4puZ
uJHlRgmTiAweEUrjM5v7/E153rE9zGQpo51fntGH5OdbWrCiPeT5UzdNp9gOiLjMtixDLI5ydYGn
hRfxz920GkqM77pNTdAqeJOgac3rMt5ghsOTv0NTwxLTP0nmtx2Yga92BSAyJbK4POLZVuWQ2zYW
yRTNPdJSrojiJHAPwkgafBZwoaQaUBNYl3HG610CzY1QIyTnU5pL1F++lx63Ng1wwTtmQ4LRfjQD
PMsBBsRuXfM7IPOuN1hxviTDz3ceFVWKTYP7UAB6Cjj0974q4sxCkhdl1GPbgLBTpE3bjspnDTRp
rU59XnPGeXQncP1/s9/D+b9/yWS4ndJfk0MQgzQmPLRPOBVgk/iXpSeAqIXsmbs/JQ0aacox0cZq
ca1AGXZGtYlAJ61c0nJUMS7MNeGz/zuLNNkRprbnNOx+MzZgFsSs3W141HQORA0q0tFluAfQZQxo
z0lkoYqVydwPBl0SkcZ6RnYWho7CKvrY/6b0qSPaYO5FKWw1U/ttiz6LK3i4CUqnufdMnkSjrX0U
S/Fh96tqz5Hmmiej1tdWGXFrQmI5g0zA5Q+O3aFqN/fvC+Ed045BdEHyUWufXO3CysD7WkVY530J
+A7Vh0FuaQWUV9GkeqEqobzIpADeaU7R9e/5zZS3wZovq1PHF0UEQoPFhKVEja7pTl4qzWUQ5U/B
hpPxGIXqru4yIFVAxdK6X3KYqrJeNi2eTK/p8bJarKhRsxQRbX3fuy0Uv3xvxyNg1CsvVqmcfMeg
qQoqSinaTqvOwrgVvT1F15zsV71mvNFCUVBhpU9YxRYN7JRc7+5Bqbmq5CX6FaNa++9JUASfTkiy
PDcXF4lCp414p1+7iBp8cbwV62AdcanNFKpJ+gn0btb2Uqj4MsdsWuahbbINXJCG8JT6K89xhxEf
kVZ7RTnlBMEgoG0jgBPFzreuHU6mGNi1DTZE2yi9nhkHHhqCb9bHqcZrZACe0jo8MAxfNre1C6X4
6NaSv757GmCBTvhtJes+KLp7ImmLOsVo3HyRxsgfcgSmDS83y/OAj5DK7szES4FZNLUF6q2QXFCI
LG8QcFn04LoOVPI3FdkAghbMNI72MAmJTl3SLJIOY1J0eGyvO3fszKhB4d5BHQP0wUxQ6SyEVdZb
gFLjUM6kFjh48c3guEPiwbD5shDExdyvtTLYW8IUQ3RrAN7wyMYrTNZKlVHcsgwQ2B8Rrq8F2qFc
ozNLwEnwFRImGFGmmGkv0XDioxyX4F/IyC3Gwu/+yXLL/4zysI1VRD1xXVLWuaeVepmMx9fLNvYx
iVoCBXQmzMuI6yFHIOTTPv3b5D4fJa8hMNA1Xmiy+svlr9JB0F6L65zM/aF/9OIc3x3bwDV0wtJW
9CLAh615O2QHfzI+vwNJL6VomShbyL7GRNKvNZ72x9q8S11LwvHJOe1IZjQShkFH2Z81IckL4kQ8
vEpYA521AGu5juCNAslPtRq36b9TG6QQX1JouVV646zcNYX3nOFyFaarVPwLvG7MviGAD1mGHwTw
vBggi33FYjB9W2GHlWzz2SMMkdBZ88/6Ci+7b/x2EUyEz2jh1BgSAI2Gn1fqx7mze9UV93pmhQ9y
DfxwhFTg7yMsnKhe8dPWcGAdS8aE5t8uGp9/09Go4QQSPOFfO1GhyhFPOYYrsJeLmh9hCztaTvOq
VOtkAKUMASXvxT3IL18CyH1TeH6+0UTt1lI7C7QLqPJ0AV/hPJPlfbiNZFS/cZ98GpmfnxQujqyE
PQBDbJvJ/UBOPt10WQzhI+/dkuxBhahwjiIjR8xkJAGMsLMueZ8YwIxTH30EOgohYQGcevGEwjen
bujjIItN+l4FHltmsE7QxV5+WT0OxzWYwxr/Q+JHALfBF5GG7SjgXTU/ITWEQ/Nzk/iPi5ye5zbd
M85RGLRx5Y78rQMj9lWDnbCQXmuEZE03qr4mhkHvhCc+1qtUqxzsn4II7T5QVu2h4i0h9RK/Kgb4
RmzlOyMci1qS/852jwGtI83+9dZW7cUoDTesX5sarDAmpoj/1YlAkqUNT5NAWYzt0hBj5AWxckW0
OpNBXyNzihcrY08lqgXDyqFNflzM/aTUCpJUc5IsustdVKajgRtivasvhKI5REJA/Kw+PnLuuW65
5hdSXJBT9LdwqWFhlu0GNmRzTzLfQLVuEeVwUWMwDOz71PueghjuY0dkn4s1arVLWBlsnQhu3yZB
9aGMFoQspbjG8DDDyktox7jDJrjvSH2quG8/c/RChxNY5jLAo2Lyo+meeNxU+0kZaSsjKPISmyd0
mEQNd4bL/jFEw9OKivD/aSnc2IR0/Rh7HmHEXkGHakEbf7c2JHSUSjokjqRWlMSo8Jmq5S5mIBzP
HcmcMiYxySNgf/x7+ip1+ilM+rjf4AEQ9ncMJ3ey9DA44BpFThODDcLWPyNrvAWtEL9WWIltKsnt
doXDyrfi8kbObhBD/JoEHsfbHZ34yzKNx8ca2/7/r02gRZRVirZ+h1DBSdEIqrR+v5nkZSMVB10f
3L8AUJuLnXaxV6G4gLnnuXrMF1Ip6iO+CmBx7fmRNcdh7vcR+EKRG2NqtVFI4P3ta3/CeoPjgkHi
tzojuFo/7dO1DI71eXGafATl9gEhuhtz6G/Whvc67gQlJzVP7V0MKrjGNYr92C8AVy+8m4/7Q3L0
IYcbiKd1rjb4HGDIIAnHewvox47bLDYdF1fDQXhMp/b+Bgnb8tAWL6VClcSPZLOgQRSCsa2WJyhH
qacFJwWkhCaz4/hjhZe/sa2DLU8moslIRrz2DL4tZCO7TDuoW3YsNNHn4B4K/2rOC/2IMtAY8ni6
N8YN7X/FUPJBsVxrAJzr56TwqmPCwKx2bF6+QhnAJBVwtEzT0x8jgzVpyJtfIGZQHMcEHkPW/FkZ
PSVjmvDOOyt90ZsvX4P/A8JrLvOPg88/aXwJe90J6fbvjxL4Nha8O9WrtHDYMTcZmV7UefefTlVS
OYA2TSMuVRXYRyiVSJUcj0N8jaRlIcjig+P7KUq7LqFu9VrnMw6uHbzMOgbnvXWo/x7JBMH723jm
bM/GV8XqQtF91Xrx3nKbjyb4kgKUlDf/5TcEKqWVti4Zt5Bf6nEZ8Bnd5ZttROHY0Scj7CRLFF/o
mvMxawC7GjxgzJdCdjqqHzxkilcNELg3FoJRppUGCxT8dp6AI0wT8dy/6UeIiyrukuFKCrU8PkHq
6lcG2KHwh581C+kUe0NQyFkyCeyJ5U5lXCZfOZJu0nFIuXBqQ26Wh1GsiEGfKE7/74i4p3Q3pzXF
lfNA2ubMRGGPtMu2CBamRSo4Y9QHeoRajTf3iL0OAJAlDp/SxlQyIDisatYyGu9Z2z7DUQkXXld3
zt/gp0E0UgBpvVUZYWsl7WUwW+n4v79+VNBiuYiTBki1l9cHIkxdA7Q1SepWCOGbfaEQotJ9KKkm
9Uf5KsY2VJDSZ+dJYBbyk3ZXD8/yp+gOXFHMVGfKmmq43x+AsboTenWAvQQDlQ6VC0/W0XOhvUFI
Xe+DXvE4cgYgNSXvWLOlbjIiCoOBEYYQMvo5UIV6OI9d13HVJWWi/EepcLofkMyzUkiH/muSk2sE
brZ91LaUBPdSIrpRWGxvA9Z5mWpp05NX0uSyfheVEk2lYoqI9za6tiWZZQEbMqAb4kxtqER38jd6
cfOHMRxtQd3W8UtMt2poc26mQYE3JT8r4/1FU7lL9lNGl1Dfb6vJ4fNf8DrCb6gHMe/PkDvahZHd
mn5oMLT5zlvF289+blLILZeu9PokK44o826KNgfkmrLzY6DuvZdchBWYfkt3gHtFz2PqUspxiPpB
VSvRqGQNnwiuW6o1y5KdZH3w2DmQ0HtwtzRYH/FDkM0CkRcLEJYNCzLZ1mdvklQybnmCqgm2nCDH
ORE4s6J50dputMcv8NfsAXwF59Rynj5ZSPrRdBtp3txXlZ0m+FBsUupoUAw7VKs1gKFVFq5XmMtk
fiRoiiD0d04FDfrgu+vFNPg/wJTB+VgbfdtukONx4Xz+sKwZLHr88sBgqyoiJn4dnBaGgMvVZLJl
/QM0tw2a0bcwXKHt1J6zJ4LuLRX+B72M4QCulTzwIB/vrdwhI1WRbIqhzQ0W/hBJauyfM2DSpflR
WNmabJHAkBMT7eEWFE5QfsmHnBqg51PddT20il58s+dz1KbiOfJ50PGcJiu4Rr61f9tGVy/wSi6c
a0MpxwjisI29VRgAmpM39UB0BnMaEQIjzrWkSb8t+CRYUuee06Q1+ADyOvcvUsepBYWSlXONwhJH
h8OSrXWlOGAUA38Ok6JNTRFjy7wbxmLP00P1C8FO3Ck4u7MLjoABNR5OBw/ol9aemboQLnrw4oNQ
eF7VvftIB7ZoUeUiry+YIVwyrApLQs962Wxwb/C7fovSGQPrdmR2N5/W9h0LoDu0NGzchGvVqx5y
BmnlwXkqBA6aUyV2Lsf+MqmVO7rUPRZYmsHp59CBxiHp3mGkrTLQDOSykrwIZ+VsePzG4dbmccDo
HtRiSpqzDXyMeh47ajdrg/Uy3D3ecHnvK3s1RBTot3Wf5prG2gpf36/O20cRJ0TvVGwUtC3oM6KO
JKIHQtWErM54QaAqt8LgYUiiQ/kLt9zQsdKdjC5nW5etRtv3SanKX+7l/l5ULqCf8Mv+KRlDMwKy
7KuocMD6p5jpX/RoFF50UbSkGV7tQLdIjwHUfMrv40jMtvxM2SPoR29GmiTnFao5hiK4LIx4VXoO
sxQZvO/KDwLwShpuyuhvyEbPppd2/EkEkMmm7WvOwpCOGBESD9UBFA98qUUL+tOm7UbKkR67XRYT
1C7AGqQrW7UVT9ILdROLNsKrNv0uP+pZ2uFERFC3oigG8V5AeD0jq4L6iqOOT6vnLuRVjHkyVama
usRJcS1fbnCbaOxglzNcOLS3G6rBpG+x0lTxAY2xW//eNQWibB68fv1xM6gcuhh0GaT9x1lpfK3h
teWpyW/xeebm5+nTlXpjMgjqWBz/FQDfUvzxIipLI/j4xmsQ7XEbbZtZHe4En0ev0qj6JNEzs+8H
4JVnmvNYosHZNfxS5DOqadOE/BtHQV8xTBYiEjCOYNLY4DpMVd4aggivojsMVT90bMCBwAgk9z8t
+YdKlpxuH89LjHBt2NTMqE4oBbMcv6+B0poQ12dE+Ptn4iac2O8Np+1og6Px26LkwFYY+ybYDcBh
upke5I7wi34HNGaZ660QTmP1HJSNnfwt3EvOixfp/IhbCpwDL1CAdal3offG2PjcRmwsasNAD3w9
Fe7DBR/12QEPB2jYWFaNgxVenUMSYmKK+uhw/0aYLGqTEXM9ji2WTTZYD6GtwZN3rw/+YWVmLJxV
QLqWY5OCPWp/fDlKd4uQO3M63Db30lVrOIRCzrtaajN4wujqQyZbK4SkyT82ITXUGvbugem2snBE
CL2qyt2j3jFzbeNH7qu1tWSVMe15OC3mQbN0pnD5DXQSv2hziNuil/G26UCLAI6wHCesuwjBlJUf
OEn9+6UxnVUaMker7D/qvgNpSGrvMs1KajaMYHFNX8X6kN+MAnhmLLSZ+a+zszETNIElhuA7Vw2E
aUeB6YiIH5MrdAMhzZp+9rDlbqC4JVtgQxdyaxx7+CwND+rzgjGtwiwHKMgCcc1s+BX8UufoU1/u
S0I4j9isy+JgdiSfbnyBSivND10/M/QuUYc6qJseDEaXneEa175SaATwEQbOzqxP9yr08ibHLe0b
jOLHFUrz8E0eUXLv7Sxd0itMHOwAiDtYdwkBPSx0vShvsf/u1Lpn2S8wXO4hBEuHj3HM6wOhXtqr
5SWYljFG1qzZZ9zvidpz5N/6moZ7hU5yz9Sig05uYKHR7UzUbdCDk0qxe/iafs5KeVTWJnAs2X9Y
XaJflmFKJJTsAxAZRP7lMz+FmXeEdHPiKvg7STSS/DgUd7FhSaKmvwRaXKfWMJX+MLl0tvfo4DcH
uEK7gmAkeUdBeZvSaRIxRLlR9ne2u6y3Du10A7tVmBpgPej0mvcVBMS0V7pH+esNDvNMTWavyFbi
0Paw7qwCIC2943yZKnlPY6imxXmXQ/FM56tTcLLlNEbNS9lTQYAP/sTAncj7L+Cy6n6OyMXsKNiC
OqeHoSFjAOT4sYJp8Gmm3MVVDZQwkxWMaDefMwGrhu7sNzaxtnKhGK9xxD7yj1YzsysWhZJYhyks
9Qdel5kJGZnjPdBH1+auAIJKWZ1OdtMt4bqZRQwlAWG2uMMZ7Ii1LCUk5oVtPuQlhbTQgti5zMpV
shOQwTFRjo2vet4UegShY3kvMqlWQ5w+ePXUASmZ3RNRtQYZnN6jTAuIRgwoYmlVN+8xFu0e9Lp+
jK5ASBeObngeFYmNjJzRBrhInKWURlK6N/D/cVEiHHNKN2Hm+NUsmh9/rHbPeYAB9R3vGvOvcnmI
bjwMOcSum+kR++FsYFhauXhu7Pxi5rbSjphjRf+9L/nYgNVIeOV0TZz9PXuh7xtZ3O2tc95+9nti
G0dwU2rwShc2LwBMDvhHrfsNYSlZ3M9WjdYXNDGP1qaq2NXulinQ0js1AVlDmPgZeRf4U0Qv0SLJ
f7ThDyen42UpUS55NrDPeRyfmPDyEV98gmzM3zUgriOCAedqkEYrp8myx9dMcHHvxwUACH4hp8nL
q4gF5+xgCYnIWlrT/7GdFUsI4RIs98Pd4vMNQ69obCIYzVkHA7dvJXB60wWlCqcGpXAHaY8RTpxX
zET+qZXe9kaVkntSa5vWEcL8AcMCPhMCO6z7TuDlVKqNpDZc6ANpOsTZ/Bchi+bsIaK8tPcfMT2g
PPDVmRSoiQ7qtZu+TW2S73CPSiEUNSQPtHa7c04OQl13+NGSylpQwwNC5+JCq64iNCC0e61mud2l
M3rNVvYRRu5Apz/0a7muwe1hKoeq4JV0SgSopSntcSf+fBkbkGJkhSL3hJMxqf3/qljPnTKnltlR
O9La6avhcbQ2Q7TEB9YtDSHhbWrMgvIwaKEON+u056j7/SK1F7h9BLAy/ks6ZkQ1kkGTpHvPPrb4
vkx4Tr4cTDGFiitSiTdk73jiue3jJ2gluyfgUpgJ4rtBp/XHtfyqh4kTYTjgJ7rYAOB9vQnwlW4m
p7IecUwDNhJvyO4OcukUjvrq/eU/Rpm391ZcZqRigdfj0pl8R3DL54hkQu46Usypb8/V3wKIi799
w+G8014IU9OjLnm8Ou4QKe3LTaN6CwhAGr+z+i6MkNTEj7wcTD1XUJDUo708L/4Nzk5piSETkQH7
/7J70dujwhA6X796jP1WvJA8KXN24fIg/hRFxPkxfevcKNbRoTwuWgyFRRzwv2C7KDsT6pQKoPrb
Gnj6WeoVvq7MlJtUuQ8MHMXG/dXsgJJYgAHPSQalmhCn3X5fIs2cppIR5quKn7Nr34O5MQ/ggjHN
qnpuP51H/pXEQczF2WN6iDb67d2yutnBCioDGCacfQQKJ0XrFSBUlHOzG9MJYyBxMSUGgRn3DKLF
ikT6Vs9glunSk80w+dBD7ZSRpU1gwDYh1kDFtq8OrUGVYGjcWq40m+LprtDLY4mmQPIv21eZ6HCA
CT6rKQKZ5ANQYeseuepsKZk1P7TCIik1Gtg2RGhLiW+/bIHzajmJ6u3W+ujkQFAOW7SpaMT5++91
GR2vukWIwwMFm3aWDz6HqwB/3Gw5CUaaYph/PYjsEY4+Dr2SgsBvyqMSSNIS60w6u4ZYKWjzQv+i
YgL5otwGuHaajAKdGareLJcZSIAs1pd+ioDaB5EKKukc7aZSTshD1Zg08+f2Zn+vh+pR2VuczEUy
exghXwPVKBQgsyZwEDEiZV9l5mqfypjt2KwTjKs1DqfJn5AuJQcBPbDGT/9ZYyqkS7HM/dEbV1LT
N3a+GtGCsJqXJxNUQuVWosIZ7/odXZqYQcCP0ut03StyqCTegVJz4HR7nMm2ulhrdnQjZLzZ+Y6e
L16mPEhDSbf5G9sfYO2VBeMmzZBN01eKZbHiUpbnNasqN7d4WBOpt70bxWEHps3Sz2AM7/m6xjmh
N21hE0a49eVuY4bxHn0dh3KVGw4BNpievZqYvspP6FfKEQRawtJ3zB6xHFbVbDEeqWCYyth0vA4g
FwjirCMEbJ0hxTwvFveo9kFMOwNQk1ye579CumbAQy0XfeLG7NJnyJ1rwlBX3qOykJ54Vk5ZAs28
zxJctiygwwrvvQZ/k1N4XI2Z+2TSuT+2ftLAT66hutiq0qIpuLazKtsrlupi2eisYz5S0hPKrlg2
wtykfXvCT3M5650XoBDQwGxf4ylzBrs8wrhurTDcRLbGiW+sRkoeWDB5RIvrwG3Umr7YnIBx+b8d
REH2cz2SuQp8fac3Q5nbBYj2RTK8gu4Ob2nVs/YeLRDZYCD2GmZZnGmD+Fl42Px50cyyBbhiI0K9
Yw5Nly9YN6RrkuHf0qDHqRo7HTJI2bzeJ48AofKDN1HrpGWLhuY3/3yW9o27I+tQhAYUkH00NpXj
9ds3U1eZu9fD/pKNKCAurE6w/6K5TRQX0AkbnEcxdT37Ffon6IyCsmIqZfZRiv+FAN86aDbWT9an
7mDbHE4xs1fizJPglt+/H3pnh4nMuBBEf/90G5ZKgJDC26fv1gUVEvq+/vaiPJCefA9tCchwcGIc
0Zzh131AAKP8vEw8hclVMTEQ4RETSe5YSwivPYzlosds9ycerAo4fcAWQIe7fG6Szt0dKnGMh5r2
rhs0zhVeYIcWugNrcqnJ802egaRJVDx1gDwkmFL45+zu25D5Zl8EHOXB3pbtej/sag0KaYCiKTIw
chKnKt7zPDQnRYcMSa5//tf3lYoMGX4yo353nDJTP55eB0dNeKIfuzHS+QwCIHEVL8X1mcDzM+e7
uebwVRESr0hlv1Jbzd8n8Dgx9FSWmdNlSCR9n9W152efDeZFDX7xg52th3Qs+YbVsO4lK5LmDeGj
ckYYVMVfdAHiHZWK0lOQUEjmflfC0d0/rMvC5mgd6chYVEneZQHWJXN+aFpmSV3qZsTD5WQRBSVd
be+sPoCoZSb6rJfGyUW9CA8GXMTCrGczNgAHOwOuUc6X3b0XAjIXcPS1T0cPa/72tx2KyL4zzoCp
gKdOsgaWDLTdv7mIUAN44KLOr6FeYJ+WA0pHE2oIl4EectRoSGJtGV3Qj14nt69D/EwMNc0Pg2N+
DBmkgo95rOLqrvBc9ZV4MRMDosoBbKADJgPYTuMnzuV3275JtkvKmtwFim5zbmyKoJ2oGrmjM1Bs
4FeP5UvmwYb6EJaxqNvdE6ByG5ceyTmWHvQTlVKynpPluunc3vykRglSClGLkAfbHPHkNRCF71IJ
c6DDmxbuGiHWq4w9ZSDcZqrzTGLRhl/GJRBqrmXy5cYS5kYXVg6wBOOoE5mudkUkeziPgdzpJDlE
fa2PJDcM/Pf524NwFoBOjWJF+bwj8lA9tCxyYmUKoP2m6lMH/TsOtdhvTe3pVyiX8ELgYbmX/4Xh
SR2NsqQEC7fgOSpAA6I7HZGAQylGj5s6clxdCiWdsp5gTQ1NAs2xHyN15IjGqETOhIh5C/fWGQTg
HY167lp8tt1uRJEsZk4U6mjNi7O5cJGAJJm8utu+L1J0QLkMR8dGlUhn1NqiLVVeRBAdu8VJJyT6
/UUclmiTIIqfKHWEBXksUv5g1DhbOLoqNtU0skrChtjfgiSXBHNq85spJwIPrP99p9EdjAYgHK/h
lUjr77Io8AxcIcS7lb4Qcxn5EVIxX7Vl3H4Xjvc05LegXYjmvwmT5lwX9df6KS+hZFGzynwvJpGW
aoKwkEJcaHim+YyY8ZL9cvaJkFajSOKRpWqodnjOUqBomJMv/YPx0YFrnVwSqzLhmwuGgwLJcO3d
A43+3NLJqcKt7RMPmIqB8wtsqwyTOKsT++YNEAeVIpVUGKp06QKGOR3gt2fgorDPKksEM/5MJ1ZZ
3ZDfRklvmrW2VQO7v5t4bJiXHK5gapfKDJBHspH4AA22Q+Cu6R/DU6b+DwwYqOWRzP0ZH0+7dmrY
Ny7LpfSOJMcKbArHbWscs5aU6GwoL9mPMqeK1QX9COBUbKgHmssmCel5Eo/Ij45FmGhnIoxeiQ5f
Bx0Eoeys8PACF5dDvK+sf2kYffDgurJCFirmNxklPxOG0PLX+p4xyLThu81u1lT/r08miM7T98Vn
uRzx+3yjb23qjfmyGUQVcCeO/tTRo7SSdHACvwhkkd/biSBisYoSuUMwGG37lL17k+1+BMY0Ly4R
Y+acudjjOHpj583MmSNXBeooLtspLH07IW2iTrWU/4EnJ1Da5FCH6QtrBuqK6bZg/igOHGUwV4DZ
ccaih3WF/61rh1EXbNRD3XgPKb7d0yC8yMEIskiYTba2l/Bg2/MglgmlKZr/VKkW/0WPF5c6zp/H
4bnNpfIeVWz+2xq9UvFrOOYv1XYPncYG2V5gPEYuVUGHzb0qmZKZdAhR9OreOlTFiRVhJn7Ad7QU
S62ZpE16s11rFXj8OdPoPwq26I4UhTUbjVszwOfHGb0ugvpsvKAgLHRHBG8sQEzHUVYTQ19/TvoT
X4D7K40oJpVm/+PsQxkIAqX6L42SB/xQIU6R563AqgbPF16HLbLdTZ56CTKvl5RUMab1S49lqSbC
2BSYxxOu5/CpcgGU7K8jBMlrAux/xIHXh7vzPC7DEtl9OET08hu6q8T3BwO5mN2aH07CYey+q7wz
OtX/mUJxacOOaXdRxlyk6SGk9OPaN+K51YlcZjEzLMqsjlK2eXzMo8OoTTTIdecny/bGO1NtwGEm
MkbScHbzQFdfrS4+ODIDkzJ3ydW0bauffnRe2+oQJp5sK79+dDOfn0VdOI3H/38cBJFTmvUJauiF
nZP+sCO22VRT341aIUfH5vVrt/Mn10wOixbjqo6RaTZK5ds1CU9Mhqe3ruIisFbz6jqZuoEjwTX9
jYAAvYC9/Wis0r4X/JwDB62CcGXgpdlWYI/lxcLZ9aDgm2k522YetFkk2ZDnN36wpv6roDbvJQgj
ZBFONu3Mep87NV93IGghSTxsFKFCZE8V3QEPN/tHXcXCWfHmWJmUNTviv3n9/0S4pNZI1pYIm8uL
1GYuKgvKTYtIH3uQEKrUQdw1x5Y/KPnoZj++PbKAFQ+M2AWVd43Mldate0+Y9gzitk2tKENCZh3W
+a5qIyHEWAhTlFmm1Q5uOJ7d0d0Mfd8np7goF3QwQo9vhP1eCprTeLdmCN66Zpyg98amzHVRKAwI
fLFjtQzlb6pGAvp9I3eXyzEShmBZjKcYR1Pg4B1mq8XQIuZGLesGE0jW2Oxq/ks35sq0PQsPgfIb
rlv6D+rVdbGboRFaMIK1Wk3aIjPofW5ejgug7apatTr7sVwTIPlrhV5EElkHem3lWkITBE2faWAg
/wMHSFeXGnD4F8HDFUXvnYuIACeTGLEqX5voKnptALA2pTLe6wgRY7zSsenL6dKyqA1nBfrtkIwV
ooKjWM/TiMX/FvEWqQwDOtJfnppKiTk7/XfNet6qDlMAADcAMDwzyByiQWJgDJFTwLO1SjXB8I4O
oYwbrlCXYG3SDvjlEyp4yi+1K64FV9roh8CgH1YBu+U9K7IaUmru0LV1sKOvtMbajsp4Dt4+EAG6
gcTtbqJnILvUMrIxnt+q9JJiOw8XW7vf2QuB/gDDlAT1NwBAcKchuyubw58gktZtK7vk13CvfjQK
UD5JjSur+99Gl+XRZ0CWTTaNlGenRq8eXr926iX4TtrKDYr2cg2wkdFrxTBsG3IS+LvjmHJyuYyv
Ox6J6GeIiXwkQkiuOq78HLJ75jpZ9V9KosQWczXo+kFg6xPc6hiAi+BMRTbjXN4vlyAsunCzJ1DF
NA/+Faw7zmUvMvSzt41TGDbzUuAvOxOPy7Jf2hccxmIdHXEhg5L+pfHEv/W8sFYz0EvbKTu6UNTA
6uylje6HPdbhBCNb11glEm6i+U3wGDRPuyhwIMMpdamttGgLFVDZvu+g7mOPlW8deiujrKEhL7Uv
TJeU7rUrbE1mbA46eJmBXF+voiXS66DPM3Y0H54tS1vxkzmcQZPHSTxiv4Kq0okDEbhokKH9kUNU
xlFuC/0eDZPv5kFBV/aQaPoxXcUoC1Stl05lHoVWgWP/N3uD3BI2AWhZBxeY1tI14PxdyEWQKOOq
mKcoOYoHJQ4wshycWUaJGLD1Zzrtzx+vlVsFSXB8Z/roHCW8rYDqRDjvjphONJlt9HmCuFY29XkT
J6Z15EN918kaB6GB8UyPzv1f3KEMEZSZ2yqcAToxjUBNiij7JRTQWGgilZQVsCWV8jG1DEotZeQF
YxkbrzNiUCM/U4Fn+iGFGpaB1QUU4JQGdjYLxSCAYsDh3Hsj+cJajz3HNuhVG3N7a9ydgUkJd4SW
2G2EiYVvkSDdp6jxNVJIaUrC2Od0ec99UDL2KxZ/5WLSE/13u91mkvJ+xJJHwpVpC14jMZLvYKjk
5g1YZQSURirCXc+sYn/8xo54JGKr8j+nl7QEh2DnWLIHbCTjjZ0BhwPPa7YoLiSjhlYiO56q1vpF
NO38bBcqZQQbtmmytW6v3pKhJ9Y4aYP+0lJbd0XdUf2BwCEo5TmiN7vMiwLdBrNc2+6G++Km/ZOT
yrCtvIxIU3qCcJkdBoWgTU/ILDHkuW4SQINb/rEWgQsGBy5AxLZOZtWMT/n2ErKDw1jZ2vacJ4hv
Zn+IdCupGlGDXpsYkPCB31mhTffB9MeMWKGLGsf3JaRB0Trc5g0odyFQCtlpn2fUj9PhaOhvBgsg
cAQ+PQUr1oUyBOQxq6HPrqEkg0tLO++O997cqocXsdMs1mNXExCNJ0CALp1oz6vehq9loPCHLgeJ
89gSiglBDKg3pXqokvoFM/wNZyr8CcI7GEKUxrz6A4BHxUcuHQmFUuue65gmNBr41luHvtKBxtcy
9SEcXsAgYfQd45FL/5hxS8RJ9Q7Hn5CRj9kiD6DNjl3KpuDt/4LTcZtK7cGsATMRVDo6VHDrLWBM
eUAnDyvvsdQrHBo+MT323B+70SzbWqT6IhlGGxd/yvgGzFKnySfSmUuxfRbFiCOQjo0SHRmpMbOb
3+XgTAJDFzs0ZqkbjZLlx/CSLdW2xVQjqsMTj/vXKy2234eZXf44wO2q3tU5dl/mbZxICnreBK7n
9gHOSja2OIIjWeG6x87zQV3jE+8EpvWdqSRE6N7/lPPmh+6LQnxf/StckaNXhcCdHL1e6KVyHICe
hz5M+Evwo+M5uXDlU1dwCPy7vjIfVusEzv9CYjln59bY4kE6XDMuDiM153hfAjuVDYd5Aqw1l+kf
5/W5ITTtGwdp+NXI5Xm1UDXrckXrnewE4OsLPDwEEIhQCH0WXuBGbUC/kpfnxg5zUW9WkgZFWHRE
xZTt8Y3kbifQCEz86HwMOunEsvx9x7cdnKDRDrDpNQdZvnUZKwxkjO2PSOVRCEtnrVENcSrjdk0y
aOez397XVLCrDrkTZQmzp9c6goDtcJBlT45gkficVYCwjBjgtP0fBGaCOieyNJbubdk0nk9uzeOZ
0Xy2RxiqzEWXQAwENyjY+JxETCxxk4B2QY0+D4i1F7owWobjASGGwyRYWv4ChsJbEZT38FeRFPfI
klRzFs40iIYjhQ+1oRp1/riM8R6pOFhYLWIrElIcqVqYJYvnEkRt9m/e3/fDpanudj8sIzEHpaIA
OnHAj5/kkuNqFg+d66T6DNbcWjBXzTYrDusXvCUbTh7lXm3CR0uiQmqQb0haqftoy6rVDcKgt/Ho
Dh1DGPbGeXUitJRWz7eh4vVaQf2WQ00CMvqBcUYVb5hGlG4tXTM1lAdO32iyRSdNR8fGjAdSkYZG
cBVIuVIjmOqWlHj+LZ2L9CXnBdiusCPV8USil1RaKPU1i69nXk4xOW9m1sJn9o8ra/rNaqymC0Wj
PWbgfSNK7LW+PNtFIJ5XzXYw6DMfuV0FqunX5gDHvRBHYxT5LbxaIpwCWArelESy7iO0MX3jxSvo
rygvmvcPsEiOqn2O7t19ncUuiJ6cYyhAx1ygdfsde1xNvP2radZJo+XKDUF8Z8bI5Q1GXfjhmGp4
qjrV6y0PbeGpLtfh2+NZptGsd3mdrR+PHS154HeRl9kRLRbxw0trf3/gLbGpvECYv+Maf2cJb7rI
XWVVN0zmdJtBzBiYXhxnFhRn0COspjv4qO2+JSXXlNucVJhuENXnX/ZIL73sSfzKvx3MwTY/yurI
Lig78PZoa5VPv130lUKWBar9d37lkkRJ1UAlv3X9vtdm/H5NMvUn71CIOZJWHdVvPAhVepOV1r41
SP02AYDvMhO1UFC0ByDIbG2XI389paTWqUMz0WSB9xnbucuZDnz8PwZdbjyJX5N+zgPo73PSaqmw
UnI9bBdM/QdSVGFqAWkMSnUUWfdlFKZyH65CHdO5v7Iewq3dNYUsbXDy8i3Ac1hKYgGLMT2zrsTc
DXSEf+j73RRHkyv6vjxIdrULV72ou1DG+30hb15cmlY2nuxzO06rMgi/w8aDT9UhVS/ZDlLZkKFD
qrnrZ0+7IyRNIJwCobj9FFfyHzKPqej47t72VBly8NH/E+7FGpPBIOVhNF44iJ01nfdr2yF1B2oD
IabmnpjCMFrXdHZyZijb4wE7qLEC/eynMV/10I8b1khmoFWY6vcpJyAq/db9a2qo/ohZxu+RCSgz
+6wsRtuuu9imgb3nTCNdPIodHVLypRpXiTPTQijQ0fTMN6mDfbGu1oTArrPNlQAao3ApZC8j3Y6r
Sp477DzHM13P6QeVFtSNiOYGhH/nKE3Ru0Ale62MClvdJJX7XgNFvyfuqbgi6vuIPa8v09uLKfvt
ueadyMj/VtmyEeoCklWrln9tVpBzu/dq+hKqJV+dgJa+nRmnL8e2lTf5c2YJ3kMqXBKK1Q2UYYAk
z/Z4l3RGhAPagRAqgeZ1u/ntlXcKx/wv2gtUfmKH+9nTh86sBWc/Jsw0071+St5wgRijC81zBLI9
3Dqo1Ua4zNhRyBIi5hiONM3WAjkiP24olBkEN5+8rxMXN0T+sYYUnisya4h+73mgfNBF5Ntba0Yb
e98b9SsjykA+7EzJzsgkSLzdQ/GAYJzqBs2Cbz5Si78DIYrHzMXckolsLihPtTzj8EeW9HlPVYS4
gWiF5TnQnDNuqQLVFQXT5+NxjmEXk5F3lCAxkmXJlKdYpdEsSi0G1AVrOUV+JgoWpM3OvxtysKkL
TVMimecrh2vItj2XCck2iA7gKSMbtt9td2I+2Hnayfnl9OpkCSbyOhOwR0U97B7IELSJ7NRNKov7
aFhL5oa6+snFIqYxEvDIi4cXF1RfoetnN1KA3W2IK2rKUufqa5fsW/5oLBW8VFqYl9ppckP8PPTu
NgrZ2SFTquxSk5yN3BjVUyjHv8feGfG5lyCRR3NJPV8gRHGRstFOAtw7ubYw6TQ0XUf1dXHdhL40
LWNPo133v+GjQp743NwcoJ5wH3WIHIuM4xItzZ8/nhZdZ8eE2WAQUnbvVKm9WOD9Dia/RIAOtvol
OAveR8qCY9RnVDbO4aP5h0qwS8xv61fwNjNYUENdUAqX+mA1zBRzyRrydWmn9Iau0Ci+yqabcepl
w3tEC8QTXcvAIu4sjN593dkBxWTrq3JkcPdX3jA+dX9+WhQKayo0ufAPA7jD4flnUgTXbgD2p5kR
Tn8Qdm06EoaTr3hYVBQI26clUmPXOjsiJQJiUdPTiUyr3HlscW++m314Mt96+AqZA2o9ilGOaANH
6G2Z76yV03U3iYEcr7SDfrP/HlsssNDgT/BXodGne0nYP1Stvbf+FpROtItk9dGoYP0G6Itp6evS
E+D9DKbsWmG89Gu2NUv20kSePOjZQvWdyVpDZ/ENJk4HVG5zDF+OWuJphgz+Gv51BckUu0HrtHL+
2ykAGu7jOyrs6iOaB2RWLt7kG6S8iAvREACUkVRMurNKDJirGKvmLbRRBd8Pey2luEen5rjzIX+s
gA80fmrtdTOfSd7AOZPLjN07tz6cKgopMMlbJ52hT96Jo/qBu1Up/hlUmIq4WFFBXVdzyFcu/L5j
Dt10qOP8wOzdXeWhgp7ck/mjDpPxzcjSeGHAuUav+D6bNtmYwD68TkbwSzMKG0VZ8mC81S59fErb
KalMbA6lUOKTLCIYpQRf5ZuCX4aqJbMKjOnF3rlQRwKnanAy8OCC8McoI9Uw1AXD7EMj1a2cKhJA
4Uttwq2bYEN8sjza9GIMnBahya8Kpz5adxU2EfIAtCfE5QfBlJvdJkjYiGM6M4vTL67iiG6tfYOC
TcATT0AjHQtq94wT334vK3LcgjnX1RB8PIRLbX5KjbCq0/aU24LgImOecP/YfH6vjOoK6fOtciIE
RtI8SmvI2HHq6QzFsdVyOMklmK4NcG7IN+lMO7TFb9NipXhzB7CcsHc5l0NwS36OU7mGo6a//ydD
zGO2ew4jQjk3ET+Feg5dMaViAnI6WwxK9aUuvuqDr1iSYvNJljez6BhS6t5phPX7wvtUAfAioLk3
L0nDMsX9N+aYn+yWfD+G7/TLcb/H7pDwbJjAzaBgaEdjVs3F+i4A65ynK2Wb+Fwi1xqRxrpkv55q
DMvIVPy9ehsHGD9rRMI5JtKA7AsKuwkPp4F4T428uAG428rL6eEF91CqfTTUI8GyPLjnvZ/t65MO
9ROv7pf1+phWNHNuZQoOdxknpAkilSXtFnyaZFNYEF923sFnB36I+vpTozWQDCV9lzT4EAjL01bM
e9hTyRXWmAKG2d4JcbaWzxFnZ7yIYFFaSkwHQ0mpu5DIum9XikGQ24p4vmDyHGW89fLwds+hVeYZ
3J1RFsO/DkkJDcSMj1zPqi34UjizpVaSmca0yTRfACfvwbu/m4goy1LfHfFhC7dCpLKUuEHO+Cgz
1tltj0Plz7MtxNv1xrpvLi8D7QaStetHN9Yz2/TPl3QqVxRCh+9YHwIrjF4CLEqKPsWOpLqdt3QF
+RV/7pLcwhi0lzP/fB5xZpo7lrgk+k95KV9bVxLbzRd355gCGq3vGMyJ9V0eQeK5mt8PvQiBDYsz
9BYRfIsMeFhi6kMElFL/pUV17awqT25E0nksjA6IzrLDHpQyYeiYJktACoBrRS/lV5pgn0LPFori
XY28+Q+6tRROex6R0XzUswS3Da3sHWzFm3aefM/JZFwckeIc18zwWTLJ15p+vDCIKRsC8QDG9Cej
uHGGwz/SA7ZH+fFdp28EaEK+QoMA93ZxZ9TLxqipIrSwnx/jDXhhgr1A+S6O5QLwD9i1fmU7cJWs
J8hZP3qfYasf8HlMZjcnKyrKhGzkDi5xEvMlgccyCduAz0hTnjB3YXr/qJOV24qoM4ZsmvFb32UX
ibmo8TT4noPqiU+cH62WGKPzwSvKPoWz2TnCc+luQsw+yTnC3/UHtD3L9WIjeqq+TEMrY+8YPnPZ
BxNTJoogTvWn+kw+wqHnut8UL1ocW5r3+n66ANh4JVB/HSx1NYIoJIRgrSiR+wP7dqV1t0OYOxA8
Rwqznmcpdk9JdO5SvSULn502wyCr0lERg0x4ke78BUg5WMkbTClK91Q27JUHUcFpll/rMI2tvXiC
i6MhGvGTq5C/xz6D+tGG1YSwpSVeP1OfbWkAGaw58XPP8RoLGBzPHicyDH+a9onTwzV25O6k4md3
KYSZsywORxTM3kuEcbKbwhE/FfjMxx7p86a2kd+9DEUm0fFYW+Lkz6HQLMQIbRMy+mu/94Jzh8D+
AV2ipJYbrk/N1UzeIwRFGUJzQOXDyCbeUFDIu41Ls6jRF6RcNnrXvdUOJQRAuYmfueIticPcmqFd
DbaEHfERCd7B0s+hC154F8wp4njDHRQPTXEFAREHVIgAEL+usDbj7DtNKKrP9tB6VZQD+n3bcWOy
R3Wm60V6p1siuUzHRpNx88S9UlCbMeukmQXFzilbwT/wwwubX4jUvLx9EdbQglkLba82+gYwzSg4
8WRO9ynY1HCgoHcqfi+HPCF6oKBIdU0lovMq9gAb5zxX7O2w0z2+RTGc7p9GwvYQObBW2pKfBOFj
Xj5eRjFK38SnindkuTRvMHlPzeuolrPvZM+0HXFzIP7XdFc4Te5wY946+YtaVT/2eL+HRmxnjWkG
6NgSZJGuZXlg1NX3WF8GGjrPVGXMxLxTnJidrJ2EpnK8ciwEPR+iSWkv1qz5q9nSEKGY/TEsAdVU
Mv3A12QBEeLeHYwDVO+dGIEbf9LKvoT2PJRTJAY/w20KlnbDvaJTkZasNSk6Wr12Wm0Lv2jF/9Sd
Yim04OskmMQl6vTfpQ0EELE4qPvW2YfrG2uesw/JCj+x7a0Y6mC4nWZFvbbImNnfcBG0lPMIfkOX
Sg5+gimywnETwI+mQLQi8+3k2RRjVm9apYf33rht89fIUWwRg6LZ6yVZxg+KId4xE2rE+snJsb7R
gGD5Ng84Kla516Logurj5AbM1kLDcsUvWuVB5s0jBKY6iV/GhqFcRKiqk7Blg8ohdqPOpMiSsaWp
dfBsHeS52iS4un5B01fc3M2Ljd5Iy4YPQd/JUPFcIVleMmXnehs8kCSxMlp4wNbYFLOL0btUboI7
KurgSojqaMw2Mroz36UDtASJTPkZIMCQ+UfuYOTICJcZ57fnEqoCHwoYfnkvJ+nS133GhXq0X1f1
cCW8tQQ7Im5UjavLQWMiC8/PiCphLq78cTcxoC5oZbHUl5wE5BvTSFgyYj1JMGwKyBrT39Crqwb5
dWFsXr9KZjbaw85lchbzK7m83bUQK6IuY0hyVbR/7PVg9Mk7DacA27ejjHOu104AQ4bmIPbrNg3s
k5NKDBEvYBAMpaOOFYTsUIDTiBVcsqWqSQ/vbia0QSkysDDzB+CIIB3iMCIDImTtOJMtqXpxEXbo
d/lecWU3T/Bay2c6zk6bXcu5PeEmLEmX2WhjzAnduQBzKTolGwYYbwtCY7nfljwTqBc35s+wdpOj
fTjIcVOSY1oqcvJITp9hCYA1W7im+bRccFrja1KDBVsc0D2pRfnkPBvK4yMbp3fZxtATymUTdWps
qvrsyYA45G0+d5AkewrSfsv67LmF40jsQrikkABMTs5C1D6HDuQ1cLXa269pArDA6UtItrErC8O9
424qYbAa6pt2mwslwmaDl4Fq7doQieqSrOJJ/KbG/1Gp36zc7HKgDpv/aUVSRmBpsrqxpy5Ti8CS
BS1AmVpOsRmP3hbmkjlYPvmOef+2k2ZFGcYdul3kmH3vBUX8RciQV4NstmtbWnq/mNeMU2mNfeSR
yuNV55rgirhFh7t2fcW/FwSSdCzBmIOESyIinCgabi40dxQOXaFDeqhDwAyf6Le0bOBrwNcdYiPb
PN0KiPrrYdrNqzRvrZvS+TjS50/MSAT18QPESiU4OcSHyxzxuPguQfV7q4e/5r33Y+2y9NLIVONx
tSE6OcN+4Xovzv/7NMUY7PsGxhLjmpS5lHQSPHrj1DQ3dyIv7ALmsTMOPnkBEUb4vdqCIQd6iC9/
l03Lry67Py6qvTse41BjlYEDtfpXEfwKtgJwMbUq4PkwcouVG1dDTKeKiAB9NK69rhi0tuyNXIF2
vIl8rRRBH+kuEdS4FMqoBjsaAN7/fzZ+z5He1vtIzEPZ9KbHbPH3YvXaB2cAuqFHNFwKR+pZaqAr
v7dX2dvqhfD0jAFcdD+Rk5HISDPqKMLMi6ohgo9mo/RfES8OFahMsxxe+DToO6QYVW7ziksAmvr5
96W/1esLNBH70MCP7ARaHEGLfAqWSC0zQxuZXlyEX2nGK+t3a9WGxBGSO5f2PMqsi2HrV6oP/NN6
IBJMzsfSwZw6AoGrjzsTA8fOT4Q96M3U81tCvFl5/AbIDadYC94r5uu9nCWO4bR76inlxBCTUuyi
EXUvhCgYDNL1RjOW76jJKO13MCkEgifFYwEKzZTmUMOGLZDgh8eDDKQhpcUFwPYRWdpw5u5o2Cr+
R+bN/iIKAQpE6vccI4BqpS0yHbBO0NzXjgjFnNOotpNDhcb6QBj3YIDeEYcd52EM3rMoWv4yZ7CZ
wWwcwH5Y9qU1c5b1m0qAfx0j5QZhsepNeRKSQ6baZnaZhUPGBfEjVSpP3RFCHSlhlPpsHp6yAeI4
mi9GSPbYWt9Hg2pLEopgR1jgQAbhkf/LapkBStFRxo7j6F8ENVbXsp5I0ypRZlD5Dol6WeJDOS41
WdMuZMN2JsunPeN38O550S9ImT3vuE+WS3ECk32lDEklKqCqkDZfScELyS4jcqXbjlcNAoj6OEsQ
TWePXBGnktpfJvbORaX+5UTIircafWkA+3DEAAY+4MKaZAq2vAFqMFmJwz8hxbDznbAvoYeu4sA0
mv/oyAkcb0BqKRrmxPupH8+wrr1mYjYin1lV0xDabThid6VJW9lSW8hCrlv+PArsPWOoguabQ2Gp
UiYmvxDxCfasnMRY5dR7YmxRxHVhEl9RtF/pA7RghXM7WC/NR7MYriHVxX32/x5z0yVore5Fag+i
Pqdt+WXi0kk2DNYHGqXEdyz+FAOZ7RPrSobapOJT9tU9u180QnbshuA8SBMRHaCJWwyp5FM+zIPu
y5xDLqw+uhkZ8NPk/3n6kL5YiErlB0AzHl2sIYnkv+RXqDrBQwerXbLXwft+7PRH5vfW4gLBpR9W
rFCGfmJTdYcmr8zOpefez7ML7IBE2OXdGcMrC9kPRF67KE7z8FUWuNiDEN1VA9oDu3LnUBtb01UW
sJSzhygjAw5usJ5DjHjSKCYbSCrOoj6FIDNChuaIlmZTz+CLuAwBONDAg1sS2iY86+b+61jW8JZQ
ZktnRul1BpcH81LlxCGX3Un/2AerzswYS7WCvgikGzNGWeEARUga+K5X1tFoZnGQCfbvKjrwqceO
Y/mo5pLGBZzI6ywvuc4iBbM/d3qksQlQn7d6DHIzvP9yS+IZJ1R6IRnerDmG9vJgTLEG1Vd2+Tsq
Q7Yb2PtCi7FwKDvMO8Z6NXlU9eFyHjZxIkM3Q7tZOhJowZhY+GA9T/bikvPM6CH0GluzifCS+0B9
M1Rm4LHBAlvrU6sBJ3Mqt0Wgij6c9q93Fjn13mBQ7PFLUN1Gq+KPTXUds5Q+bCx703NUS083+x2V
R1o5pGNU19w3ZJ+lfBaAORghzVmM00NPgj6vcVTBaaoWb4KhaGY71OYWYYh0V0OGPzelb/iRQS1w
dLnPUcxKIVcZ9WWYXa1m2CvG96bIMAvJOdMjaXBbXjeOD2aG424HZh/KNhs5jLb2nzleKamC0p+1
bmglC0Kj76IK6nBFcEK/6yqOZRput787DbtIJU2rfGxfXqh+Igdj3eRPSIS7SPfXlYXEeTV3MdUF
BK+Ehe3+vj4JqIx5DMp+4UPkbxP0LiE6oXaRFSKpWTEFR2rwvV46N+IymDLqz1cJ5EAC9o54ET7S
EqeROl85kY6RD5yrwQXgcwSOxRGp8txV65umeoT8krS4+kory2EyOXtmaCSp8XaUtTMccv/MgTiT
X8eKLWm5hFuk35H41ioK+rY6RAt9O5nX7ec3Ce2sTPoLwzuXml92Olvj40GX8hZuCrLL/kWeheLe
mGnLKqllSztndI2gau0RlZQczDPZYTXwIcPxoSxTClNpBy/OGwkKne/Dc2zvDNoWMOOtYsqH0dTT
2CM6bJdYCTCGh7p9dXf9hEihteq9l2+xuTXpvPhMzBpRyuq+8tPSs1s8fFoahnJGlZ4TnybAQXZ8
D/D6ecj453xqF2AYg0FIp3/GK2sbGO57PqQ1rD3fyXcyP0WYc4xJJZA9rmwUHsSToQQum/DmMAwr
1f8KFqnq4ArpNAcNZq1UBObvxLq2O4czfhUiHhpcqJ7UW4huvOBon3ot51x27fImNfeNpBbLmFZ9
0LlxlgrofBGfEIeMe5gsyDKUMsc09jyBE2F0CIeJn9W2v/KlruY4FqH7t2K7/PFPcLLsPWb2RkAe
LMQo4Do1+M87lziRk+sNUJX20K8ArURpJEHyeyNEQsuec3EsXi/ivWW3YgqATbp+DVSN91o37OUF
9kHS1ag/Ps+NAHaGf4iQVQ5mIgd/2GVr1HrO0EQP8GZ0zHrsZwgMESlq/mpTx/fVb9J0NHMT7+pu
1wUlLU2s29KqP9+cKzFty14JD90SikZEe+It10wlXuLRl2F7j5TmL546xPTyTxwIe/Ug0yErgPDY
k/681uxD9lUbofLnT8PcwDFwn3vR8sqvlW1EglHaUFbtCLXcsUi6bDJosHpHZERcLk88TJ+ADxOG
p03Scl4tjYxTFvKoZb77Ofc3iMFj+j6XeFUBXqZc14SKxPJTSYmuA3/466kNavzJ/5EIesXqJEFP
fPz+H009qaSsD7yLPjgx85NEShl7EVFj3Oyo/e/xIePQsMUl3zrA8rbi/Q2hcO6857rqBpQ0GbWI
gH2j+kkXi9a/CjH4maXtLpIczq2x9ZChKdpPoprHFW3iRFDcK/sQOKMU/VMm4A12awEX4dcEur/i
BovKQV84FX4OJhi5nj86emULeQ11tiB8seE94/gX96i6BC2WxbGVCBMTIPMCIAKcVxmwKvDgCIYM
SuJOGQW0lAVEgOx4sFSJK/HLdiqJjH4KcKF477FoiUD5prhoGYzkeRcBXVqL+PNCHWZo90VH1K5i
wJVW+6ElBzwVCPxdVt/vBeJgOk5zYeM/uEKWxq6UB/atKpahGf4WPZGQFgZpyNl43yAFSpfk4QCK
Rv9W5ElWQPGDnrt4hT0oqRzwHpXZjaJeEzZAoKcdX+uG/pjEQQnGzEh8JBEqWgb0sL3iFLm7X1Bh
VqtIreZLwDAgT1rJmMUs65bSm8wSm+5u0lKuhPGOhP5sSVkXR4IaIzk4N3i5iJDCX6eVDxn8z6m5
PxrCILUQTTpIOy1aiaCikaAdhJ5GkFL2oEdoPtkf2Hkg+EPFDWDj5f7pUGS+SmXJJaUFIYH0klNk
PpnJQHy6wt3HgDChjWunRGjXqwhAIC50Y+fi0zU94aqCIDhwig4ES4O5vJEZjjjsTQKkQQHtRU9l
vemQD67wD0pN4wdzXBifoeGoqP5SjTgm+JOZypBVv0fn5eq6e1W1LPiwRQikm+YegWWd4sZFyGNz
Zh9hic+F+ELHR3rLOdCbzGa/vvqcHJtj22mAGCyu3iB9eVVOXuSHzck2LggLCOqiBd5RYpM5ZrqO
qoArbePnrp5fGc39yhvKvtBZcKkP5DkZhTGEKFkPtpDdaHeibTNOucacL1gk06E73FpkY9otsZb2
6MZVfZYN3L40NOxoIPgmo4nfFGHUTNO3yAMlf5a/1gqjtdqDI9rWu38LTmRHk6eXgNoTbcXveYFs
VZcBcyhkwoSGVoW7/DKohYNX1LQhZr7Wd3o8gk8PvT9NtMYO8qCNP8nZ3fr7xblC/xAn1S30dRKx
d3AMYQ4H/cE/wbj9xutEZj6ChNN+rKCzdFMoizUcfBaiFkK/0+jsAQhXKEPX3K8z7xCQRuk4Mt7G
3h6ymk/TddkHtSc/eu+Ez9ztM19jmoygMN9vUwzE+QIMfeZCyCjNl/cnYVoqcWl2lGliMMX/qaZS
CpL0/Ej0D27LOYJ3dOe1IbK733pmHGs8Uyjk6vOz3YAWiLWvqbrUmNM6UW+CyjAEej421otExDq5
T7S0TG/Yl9o3cEGe2scCgVahTibfx4Ir9+zeLhkBvBm6d91hh6xWF3YyMrEXQFhAx31PA1rHnvtT
xe5rZy8pkijC0q7V1Vsc/ZBMOl+0Xtd3ksJmd+hZCtYI6mKd/L66UqygwyEwWtrTbvxhKpjlLkkE
egcQoOAvi2a+N839xOFmhcDUOojHm1eTh0W+8yUcQWJYDarZGUTPPaTO3cZbi5TtPSRMu8uMqAsX
/kiiet5JgTiS1roco0TEoS5wmw9l1fZJHvdOYGbwDx9l/vjV4v1KpquY2aZmXpxCIcMvGBp0bPGL
F0Ho+vTboPghwp88HlbKg/dv99NQno/H2vW8hM7mcExY6iFtKrwrUJEVNrI49DHWhCOPs6LiERK8
NQaFX2QzZAj01xTpAe3WKS985EyePrh9X4/FydlZOOtZUYlDAKXX71lD/uUZsDNACeOPuxCfZka5
aNFYX39vLDlT10tztHfx13U9nZa37XsXP3bu1FU68nxHJ2JiZD0R2fufcXs68EtysNKSk+nsw5LR
FIgkgotUUjKU2/tv075Q6V9AwD1MLJC1OYhey+MDZUBCq/b1LCExGHTsolxcOvxEL2N3cFObBpc/
nC5/JiT5ejDpUsyj5boa1KySvsAAcP0CB9XuXD4TGPcjox2Bb2Tfbehe6b0dn0wS0NWzhTGRiWFS
ZWDmKbTgKEOI1VTK7+gcPo3sWKB2fBv/gNs/HKlkH3inVH1KHDkAzgfPjnjJiRcOnICkDuLCzZPC
anZbYFzZNLkZceB/9fIQnhlHLPb7hjKGg9MPkVl0esmNjKe0oHMgETuGBLlQpz66M9E38f2gCXg8
x/hzWuNPQ0or776uTUBYQH+6UnTxkRIT7jrScaNOI1rNDbty7cxf+mpTwsBzr4/wigsoWfcPTlm2
KlTwxubBKZZxfeefdOiyOjREQ4sjM6eTpRlJDAAUqjBnz7MWMqW9vVppIUvEaW74O1jwAUnTtIjc
NpOOoNQLNLiB/GljvryFht9QXqf7LYbIzzM1+y0MmTJYkzfbpONYJaY4D/uunNhBSBKaYnrSSAZ0
wTSEF3mLLmjIUPORSYmoKANtKwLPlINIybXF4V4kAdeBtLJBfk/VxK4mHieRiBbbPK6XTb8Eve8e
GfrWOlz1PxrUhekDfEkv+TXBfp0A2EH/Z5AoXTNjJlUrZwJ+VafxKa808Go1Y/lbija4TI95h49F
g7kfCqv4b6BWwivloBiDMs27AmTLEVucV1MCIflGgLT0Jc0ornfp3LdhGscfA+OCP0c7n8sQf0BL
SMEHbSuTZv0vyXT5xdHSCnm35ZNk5og33aZDjW2bgDVympjGk5rr6dYhCztZwB78qv7bFPbwHLsF
XS92IpkSzy6EYtb+sD6gYVmEJT9MO0TO27UlFlUE6dzYQPyaUpxbCG4zy539KiqPpkIlR6JpV/4n
ON/xmJJg7HOtoSt3fO8Gi3AtFDu3d+1QQyEWrNMOokmlwxxr5ZAzqwy6MKI5wUmI53v8NiNGSMvL
ppXsaEMrSkpAlsQYD9s9rxPWjiR517rVIONrtu8ifC7G4MFbsVmcB2Ypx96IU68ozFIvMODQvgrM
f8IaClsmabWA49179pzxx/3ESv7LQlK99Pqz7QEAwLJsVtNHVvQO54DHbYjG/awsgAsK3+gqQ/dK
JqJFMu1gyR8yK7jAF5Srrk0Q1a0/L26E0n6i9mrW9NQVzM5T3oXg8cEs+DA2/FOyrXq9bVJLDiNv
byuleLz0E384va6Ny/ZCfOQ/gIw9h3lp9OhtaQW2siljraur/sfxTv6zthgbqCai1It7lKlCUWz7
zGKJgbj6zW4xvjOBdKiki0mYwMXHfPsqdP7bmi7inIlKrowG1cKcxDyv8ndQkN3tLLRXAiVIuh/+
ekkYZiUOKiy3owPukgRoBcTIZvGU4sPPlNybFLOEhVwVQQhceUIhdv3ENmLvFq5CRNGa6pqdzm/f
BptaOI5Wo+bYhxWK4sVkfhgf24CUQVeyFj9TzevMJCWeEUllF6ZUYsFN7KziKbZLT+zbI0TaoTIb
fJiV91Tyy92affS0smbQPI1j3y0bgWSy00F/HJ7fOi9jKcawb9CUe5n0xaK+uXUxYSgrNkiuSYr8
u+ydovUIZLX2wRWl/Zag1I7IKAwPgiYAVE53FysswhoLc/U8erzlYNcYES68s3R728qxY067ffu8
hhSFIbAJvf6ZHCKL7Z3kAIbbu9Ks1k4vJHwWXKuC9lNORpFDVjHZTvsdPChLUiNZSWu+EyTWZmXQ
0UNmZiad1ZjzkmorXee9Q7v5JApX00a0RpmOt5AKsubThDv62tBIiSF1p1qPbXeHUQTAHNacwS3G
0hhVenBTzjF9MmjUlEGhvXNCO14U/M7TayZmv/2y3bjvpTeqkTXZeXeE79hp5VbyAFhxouClxx9V
+CVTwjo2VtPZC+i54oXXMh86rcSDou7CZR45OImYlBy9hPTBlPu/xUxzGaK8NVEof2C6bjNuoUJN
MDGlWVQe+wGi28re9LwzNEVmN86uqRPG/iTLqWvUcgnivHsa0bHuZ1eA//GnqaR1WIeNUU2x54Wa
qbMQ7vsxfmJI8S2QCNoccES5C8IqbylU4+mLbG1FdOKLSETL+8wLe/mxH7N3Zf/QIl4c24sOD9wE
ihTwnEhSEGD8TEpbSVtZKQDIm5FHYmEq3M89vOngTI2ayayUveCYtyst8IV35Xu/Sw0Zh1eNrFPK
AcileEK5SWmJKXzd3HxDq+lAYRRdjDIkJQVPxAfwIKNIrc3+UXagpNY261KGl5qvKGhp2QlEhKup
XrKKGSY6LZ6/w+EqkCFo7BSE03w0UkM4lNrIfGJTVSU2bFXi6i/Bws7UTaUyBze+VUXmqeuSqNad
HToNwfWvP8jgIxKQvWFl76YO6rISI4BkzTA9QM+7/nhb8rTO+jhNN9ueF5WO2AUMgonHKEvmyXOP
r8nwBC4S6pYX+ckBPCyYFXxBQatvOhf8Gmyp97facofiJHxIpc1WsvscNzc/+FkfjAJuAQZmNpAB
J/O+Ibr/vzyVXkFIVTQOgqtgr+26/A5+PWB6u5YeR+LknIcXbvekLML3S3tILmhxdGPM3ErDQHrL
9rbASek4IZvYbe/l0ABc9N5Q2pmBLudbONqP2O5/KtK2wMtl9fKBwVSg6YIsAQ3aUjoMC5CWmuXp
72dQJ2o54ZnKZCN6omcsnHK8p0bjn0ZZlN93RTf0bQJ71Riv3j2Af9gfUCeZm0e/O+TT7n42Oc73
tbSIkH/+/W7dansibW+LR36saX1r6Z4hwSnvC4Ge4jR+6UvmpPof+zpFh/rwLsClJZRis7Ps4puN
EBaYr0lqTNjMyCy2JMGFNHcjOl2dEet1ZRrZJEsv5A7xDNlOr+uWVFOsaWpKzYaSl+9DRG0kOA0w
1m9Slk5kPh5aMop2mqyqQDhiN/8YleQ0TJCe4RD9d2XQi80CxkzuY1S1TZH4aMs2d//vuiUyrZEN
VY4ZAr+MFUEQ7osyZcpnLMXEOv57UA5ONfFYKnoMml5ElRDb8du+RmXdieIdeIKfYjfYnySgtb/o
JPtZ1G2UqsAQHTnLyYivBZLbk8BxnypZ8QFjNXAC+wVMIxSC0Y79wS63xtsJnM4kOt74V1/ViGKK
nctJE+pTUsAMtKYBjw3YK4XCVW1PtpsHlvZ3Ce3p54YRJMqJzmh45iQTgaOwg6E6baQRf7HG+iJw
3nloFmBwhCae0RKJOf4PBMnNXA54S0CuHQpENDJMfaY7EerP/eXjXaoU//Hn0VZpzM/g5wMlfMB7
i3Vs3jjqcjqwBXXrbqCsywHxAOdQrP3qCfMV8Cl7Lo5V/KA9F8DWmW6OWRwgnBDjhKnr6YWxVhxv
7NErb0pDWoyIbYxuMAqUr87WFFPdbUROlQyAaDTm6Ca58aGh2RJMGXPykWlONjXU25+bNjrm4EJX
Qs2lY1mP+LxSoq5heC+j36boZeTC+w8rwkxBf1xvfZQ3mINMSWezwlPz5lDq/9WDun/ky1NK9D1o
rv9vQAdR6m8nMESzJwm/eNk50xszQbbAUjFJ3CuEti6WHpbH8w3RQo5WhmAR7aLMYmeJ93MkYLE1
rRN0MEz58DobLB0dTo5m6Lkkn0y4QjPi/m1qpTsnxyyGYzOjCZx+OiG9dIrAgeVpfdkIsAsN9RsQ
OzcfB102sNUF9jezXwTYGi55XU9+X+7106nXdSYgeHWCor4xr3qU9c2fnMVVoXMabt182ANluC5B
hSIZLTh0M5/o9j/ZlpUiqFSrcGdjVYumPao7pvs8eCf5H0sOral3f4t56ksm++TOw56b1abdrpU5
f+zI9ii8+t3x251EaSfQuiQorRPk2+oZiQlWpIpqpNB+YEAFmObOorjk4pMJQ0tXHcI4hyqd8B4l
bBmzglLYa3EuMKJ3ylL8woEXfzzLNw+pPHuoVaEZ0V/KHTv1Q26lIc/+4CFF/9O2ofoi7nVkNjCX
Muzc7u6gYPua+VoHJ/WR+nykFUU26stv661aAjO7+vpRENieg51/OX8ygwU6pOPkTMDvVIk2oibm
gkqN9wZgzZ3kqRRk9/qvRVX4Lks1PPdIwlm6RHOUUa22zoxMzHsY/48Eb7G2QnqNpvnQ1S5tteJk
1y0yzquW6hEtvAeZLHRgjwuTUl6nVgIZhUXaryMHD46+OcT6Q8mKvlT48gEbFtQJGFj6JX4ALb+1
9mViDavmxz/UhLRiXk+cXF1eVBa7ckQq0f5kFG9veUf+ckXkccgjVceGgvmv77D00nO5fAN7WSsy
mAhhzgWeBsdxNhWqQhrF8wruzE67JuVZNv9Yz2fKtLNaaK4XlGAzMH0tnY643z7KzgQ+ywRB7HFS
ubasWxdyZ0iLIiV+GOCIR+/rq6MdBHgQWPK3RON6gAzGyEzVFYl63DoX1Em31vNtwIn1dIvFSkuc
qa14iap0qw4r//aNzpy+6ZK3Zd21732sZHpGNaUmXA/whq+YCclaxdRhQ4+LbO6EMolOhg4Qmsg+
JORBx4U1jabjnGOm772v/yb5XrLC3ldP0kqWfeG9SoK+IcpwNQyTEKDObkb7Et0efW/TeEJCxqV8
i44eKuqvLkNNlIX9KSnW4WEC0xpA27mAmvNTY2C8eU1pJyLPfr2ut308gbsoAXy6Ummwza5vqnO1
TKjP1M+3O0yFcag81efc3Ut8Wi3K8SV/xDRkNcYET4vyj7hp9k/SmUqjNVTHBtuAn8u81jx2FHkg
LF3wNyr//f7pYpUz/uWJUi/lbtY6xzS/HVUDs2uDvx1A8bVH0UrfuOFn4/ojde0AIEBbcP/2Ux2J
Gj3olK2EYrQG6wd5WP4JiVKU1zDaeQZrCNYjMczsiWby/3X9p2q4J6yv2D1T2wB3Q73KKak9dl6m
Iewrb3l5cz+lAkygyKj1fKVP5MjsUhviNz4IB3TfWFug2H83GqosXNLSgZvmBrdwpUTFrQ2Juvj8
a+zEXMxk2qLsTPH6k5dsU2jBplVcgdZpUsVm3nkS2J3GJ4VoypChI4kMaGp0di20V/G0mQDsRk5k
zBTmFnxJZ6I6k1v7sSGfubYTZCYDcue0yGFYqjFBcapDYhQxH4J3Wwh1dEFelSECUXUXNfTm+MKC
6oo5xA7llaRxpKXOWyW3YlnjuPy2kSI/9rb9uzeCMp/sA1uhi+7OfNek3ZsBZAUTrIrlRU2KJaxb
PQoX9030ELXutE2dybkQWfMWVEd+WQabh2P2LEMcQiGbd0zIynFhU5GtasEHzOh76jhSuFYOlpVp
fSykI/lPrjPMA4P/eu4Me5B0oxR7OZHsoocE8MdYDQG1EdPSFqR8uQaRIK3cth29PfOsM/4vyUrl
yNynzOO88v1TeQTsjG3rBlsw7f4+nwz6Q6pGMPZWPJgtIBb8lCapDzVKjdMYn0z6YpESvdn2CYc7
lzCnuCm89yynz1ejs2vH2A6MnszeZsYe+xjrfxwg9rsMjPF9MbhphpKXTn0tBa/w9PAqR08fOgLB
A0EmoHybakTr2gVtnPn276CeVWbqsUK3JywWNc8YToCh7k93GrBGAsZ/RvYhBH1olsuYn15FC8Ba
COUX+ARQkXee9Zgw5FZLht1fDxN4yPzCpXWq3LJDWYVCurl0S1dfFl7hKoXz1wNQTsW+ssHmpPQV
OOM105/FFMQXkO8hfnpypEMDHtdD07GSOdF45pulQnE2hdvoK8d5JP6kfxwS0ggI+aZWbq0EM/O5
CeoUNittnN+5HVq0bRW68iWpZAkOqUv2oCOfrzncnDdXu147Mj1Jx/Axbg/CcutUsEN2A29Bih3x
c/3cTm6mTimAmcrdkFPr73dRs3w3HpIDN59FJdx50jyHGmHcBWZBm6aZY8tqGhW7iqo2yTwHsKPc
lbLnY5e1LHuP052hw4xcjWWWJyBcF4qA6nkyw8YXx1UAqoPs5zJmFqNQ/Xu2U3huHV55sdKBt0Pn
cD4ObSnUplMVsHZIP3/mORfALeP2H4Rdwh53N9w04Btk/WBcMZBIFD+pNwOYS5O7vmlWBKTcc5xX
9whBisixhrhfSyDl7J6k+345csTA06JsuyZUw9UjN1Z0GizOD99T1fm60XeKT7+oX2A+ykRfT/Jp
HYUXAfaZGOzSZ8lf4mY+2MZlKZ0aUvS4qJWoU/DAEYoc99I84NSRBYeLkmODHheMSE+n/rIZY6+H
EwHffUZkyOlCZlwiVzyx+PxALgR5+4QIuRBxnBSMIqPw45b5X+WQNbc1i+jKkHNgfKBdBryRkL1K
6ojIIZShOjgNR0LaVDbxX2/DQMbYpL5bfX8KZnf5DPjd/2iLjJMy2+Z8WqWjPE0oKvvQX/N3iNeb
+4ahGeE1mfUCu7bSeYWO611QqmwtBSG5gCMZEzOROdHpiC/ks0nH94Ih00oBTSjbK+LqvIMgCcSn
SBffZEEoU/CccG2UsPHtXaG/R8ZC0N6TwAET8zxb1iPUQYEZcOEHpWPiZxe3dD1PFHgZT0CUO82M
BaonCAt0fe09Aid1SP6xbPJifJENuLpdKXEoi4ibGbFw/f0pLICJlDK2wE3gcQa7djIQ42k2pRE5
VsrX2kI9lEzM/l6gWwI36THM27xw6d9RcwAM6YEFkFp5ym2H1ajFKp6+urB0qN5QQcfaG6iKZk6/
88m6owMhqNKPaRFO4P9XTFctpYb0qwfUqErGqPDMs454f0ff5g0YQ1lcykna9fGDthflWHlMlUkY
+yF3wKePHNtrt3/uJFfdbhQnAYAF2eBGrri9vX6SRvMKaxtlp1CvzuolWckyku7MKNxndJkinqjG
ZSdFEE+uxmjlxjkXDHPwE7vvMqqMT00VYCx8OjigXMTOUDLX7A9n0vDKfb/8oAicysP1uwP+uB+I
TpV+gtakoN67236dzU8eoUXGaQtCqEe2SLHlhW59RGMzZ4jVld0BEEZJF0Vj8daoVcmdMJWTlHlr
EeBnNt13LT/W2FOyVGXtKFfid2q9NTCQLcEbWegzxfTclxkClq+FxtGzkW12Zw6WCTTeIKBImotj
kE5cQizbdPQddVGZFNjJ5yjk4Xcwc4XTeQp79NOUAerDuCDiRO1BbOo0FOx+CdFVuhdqD1qFWjI1
sXi3gg31dOqd4J6222yGfqv1TRtmAzhodhKNdhpTi9GUNppfo7K0Qeitf91JldmojcE5MHw2n9zS
8loTXWilBGLAMwVs+sGW6cgVApfwnOorRpkB0ymfwc/P3OGlViCBixr6s5B//d4Gia2DTemWgA+0
VLR0v8+J13a9LsH5sVrquUPb+zuw/FuEHxnG0evv0zfA9w9e98ECvzDpQ5qUvLqjZEmDpKhJwty1
22PZk3ThOtx1aKV2Z/N7aali5FKQgDSR6lrKs3ljsvO5ERVy7cZeBgQgdVrtTJPqyLL5w20BgqHK
0xp0PQUnJsoaAjHj8UkRGUPwklBcSXuXntAhCRJxp+VkHLDyFERHONwx0nB5n1MiZ6oCUnI0s4ii
ATWzBw9ztZzzOQYP1j2pwiubK8cRaRL6xMvKZ8DvOnzvKUpO1fAhFQgfNWLFL8CND1GK+CG9rmsv
pzQm8flMnIAOW6logwe07cIQsBeSl1WQECEi+kw+MVeW5BTSzCq9QBHwg0SN3Fh4TfyoUAyvXVHy
sN10+YXkapxgkU7IFwxz5LIb/OuKlZKFZhNNyzqeO6j1ALHZfzHaKQYNclpF6S1zAV90tF6+YKHH
Kt9F9o5gbQAUak14qGquGD5/cXnMWP2Yj3VwJYhkB873z7QtrzHJDAV8o7r5pyfDhp6pS/l+acHm
tvB+GRzbrHHJs2AhhuefXpB2IXDkR7zUbkNgaLusC8BeIHTeovDBAlF3tuKuvRR/tyVDcgeDXnti
AU8M0TGiB6IqaM5CNUkQdMIFw0mUvf6e9BSfn9f2qkLbr+DwHaeaKMu8fgyZwBxmZwhUR9VWHblJ
lfhXcob8WiRhHi1wKMKROO8dNeLZSshfdj0Oee99AmB7YgYCSRYMD1FLQr0pZbEUjr7BYDRPDpYX
VvSNguZWF57G+4f4YYWKPxyUwZQozREVTNtcPb+LBQaAz9cA9PWNCErW1275+vSjG4o0XqsPk+Pr
J1li9PcuKcFMsY8//pj3LTBHdKEJ5s94iF95lEkEHuvl3Jiz748OVwa5gj7YcFATWqUsLAWswNvF
O3tltKDCg9KNkc3x6wXJnPkfCkOL6IffyYMU+cbaKdAhTpIX2Uoe1cxGDTJ3xvV6MiXu/wnzxrpV
DkZJZiDLq/fwXAPLY4cqnwAZa6uZ6LO/FvJZUvBavvrgBlwu5qbbyQ3RPwGLrgJ0+XxKLkVuRhx7
mNBXhEwA8dAZp/6p0RfPsg2GG37EKneDCnO/zwpud207bjAduOl0IeGSvqiBBWb8bn2TRS2tgfxo
FVvotlt6NThVBkhZrb00TWdl2Gt1YH3rbMwGKZ/+WaPwFR4f/7UVXMD64M1Kh5unUlBUV6dlUCIN
8VMku/jK7uPe6Q5GbzfXFoZhJ+cRbj2S4jxCIK80iyR4K5/jYe7g0IehwpnKbAlRmTJ8qSF+pq+g
M87Zeb6uDwAjx7A4Rv6jIPULPw1fuCvt6YGxVYC0oFRyBTiXRqU9PVbDyxnnx30HwBliMK5OsTMg
EVqrwlDN677yOout/GSELFE8iZlLErJ+djkakzl32MkdPvVD47PR6RmWzV1LAHaVjoIHfB+Roo/J
NZNbQpp4fuq0DVX8PxTsJgLH+Ws6XNKLkWPRtTZ+Va3DhlVGnOA4a/z+OarzZwZpa2PgofYVUIMk
brpIs1UixINvysqvVSUC2ljRuWsGVdE4EbmgFx0hkenEuLKnwuVhuBB7nUDXLBmcA0RLrzzOaLD1
UEFwUn/ajJ1y7ttMLs/Uj0nwmu6/aFO15CJpFwfPJjZh0lPSH3eaHA3QQt+f4OJd9uUyP5T2MGPL
Hp0dBg1AjFI3DCBEtGX5h+SvxxE4ueVhdWGEOJh2OtAviVlnd0yKkKzAsYZmcW05hOEL+DcAtxhP
f5lu1IrJFubnICgZv8C9LlWiUnJNUCg1nX0yAczvUEcXv9bRD9qfh2PCm85QqlzHpbw1rufcrYB6
9zVzyx0kl/7Q1p+zvm85Fj0oxfPEcs9HwA1EWfw3cwCdS8t6YPSEfYtA4S7xjCPfrxkbnfNPZT+A
no9aZY1ZwNsm1zQKVSfs7NdP4em+8tsU/FjljEp2haQEEzPpaLW/SI24z9uDo/Fi97UkngVM8Z9o
/Stha2n1GwAimc+lSTA9OIbrWxUwTv4Zvk9isV4Horj6VVtrjiwuTqxdp/wH+NYiqwYn1toATkvV
4C7wRHtWlRCKpWH6jFzIpPyCUZGs56OzMW/sMMNuopyFQhVOnJY7tGdPumNovQ15m31aoB4imz6J
LaJY2VBQKIaN9lZOs8Xmgw+fRQPCaWWb4FoHlVmIZgQGU9q5C8OfGLkAUlm0RNk1DHOGo/isv9xX
LOBA+BX4cBTAxXa9kagDY6/cMIaZTbOIohxyLvB14fADnQGWkV3rxy5uUkhGKnRApgd9x9/g/q+9
UD2MdyT19+Jmlav6+oH0rSsmJ+ciegSoa9NEczv5fErC5t98trNr4LmoFtLDhkk7C8eiAmPP+U99
7YBKc//xgI5Zyc1eyjXfYgYGoOiF2EEx/vAX+FmTW7Mcr8tKnIUssb+zy/2SUIroCGFSTFlrp0ku
8r+cSd2iUQddjVoiVm3yrm77gT/v5S9I9TVMrnM5SQ63dYi3BoyvvSccas2vy12PlY0dd06Vg7Eu
/SSEtz6XxzoQfTk8Krp4RIcAbT8AfgoMWe6J6Yd9L3+D2CJ905bfFLa2WhTDE/2TE5peZao8VDSO
18gXeZZhs9Wi9HICGAmbrwE5j/jU0LoeXdWHOUCTYO7TGd3MUE2q2zidNp8audjQSjW6TtiAuPVw
BSZ5hTXIKrWuLuKjU0szV3rUMoQVCtedApUUVhf2fLKw7kKyMH4QMtWgeh3/8TPI+b1RgOUHwwiG
489JU/PUR+g2Fn5hO+JTqp+8FVsInISquqMkF/ZY8jKihF9cGiYceCBPtApbdMdlLTKAJejLCAIv
IMcjo76a/Vr5lmuPvwy5YIvyclf26fyafERP8LvPP2x356DjPm+IZ9ZIAsIlqvxQ9ULrlqQrpu6w
eBsaXqi8y5N7bCl1Zj/K8c/N9BMYch02ww2BI87GQPxyBm0sidxh6rIXivhf42I+0h1QCMIEALUT
1J7SY3yOFUpGcrWg3HUDcfbee06uInvaf1kvGtmgMajcjAnAlPqmzcLW3MNAblGEQuDxuRKmQhyZ
dFMN6Pqooefx1otjNWbx5+bycIcPOEK3k18wurTcoUi9GMdH4RZQ/z20qn+qNiCgtkWQq87ictQf
RCank/0RAGJRAZY8k4Zkho9SLhPB7n4ezXHhAyGCQ9oTplL1Bc8Qcuvq34o9SOIMCWSdaIGiT2id
Z5pK/vyMvdB/5HCk5q65OAzwbiGe9I/ArvVXIaXWjdmg+Lxm3izuaRJkv1F85XVIW/Q3+PEwNEyI
SVcki+jalU4Y3Q4aKl4GiU7w2tNs4/B2C+nYR1vMpFlnU+Ji9+oF/GdKaEr6NNHazwaWxXmAIeQF
JZv7W/yodrADcgHPCfsyYRH2gc6MQm99HR8i+snkIp2fOGs+ypuUdKVf/so8a476wj7htgxinIFQ
nvi+/I6xikim8CnrpnBGH7X4vScxtfNhUGJDXu+WUbNChnssaDiQx3McG7Ilk4OFe4GGjEg1Z0g4
w0ltmn5YwvCrI8UsQi2A/yJJL9jsUE7F20qIyekkaMeOuQkwTSbFoocQ2dMyaj3NOiNmhf/qWnqN
dl7fLUqPJ5Myd/do68NN7cFJ7c2r53iLY2XPx98t3eBAJG+fQmRtPSb1bRu+rCOHCjQ5FwfZSOZt
bW3luFGXGW3X3D37PRhGDYn+ihakxVBNm2uxrrPzXKornC3pH7MnLT8gWFSdfWh4Zb8F5JH1gXRY
nmC4NSQrzT5QLSRa5NolGeTaCmIPBQWlWwPM1wRmBRSYkyCWcTUGUHTqrcj/ea3bQzW8DY68S2ZC
9NaWRin9ZJE/Ns6gKupxEWtOLdPbLlTZ6aWsxdVswQg4gZjPWiCDw6YrkE8oxc/NC27Vy7/X1MDb
H7l4/39jAFtVH+ycP7f6XpUKZncMuORSvyF/U7aLG73NVx8/DHKyT6s3aqbIGTdW3m8hF1wx2W1j
/mDOE0/ofXK55IfROjelGHEYX56jVeZGlqtSUVH5kP5prN1CiGr5j8t1IzYQojbXRbpKLx02WFsn
GRsR/eSaEe3yBxyS9SAuLajMy9GhUULhYP/nSp5a4gJMi+w0L8iShsFQAE4gMM5yDE3aGdw6XEAc
mSkBK9oE75Wf1VjE1YIetQTMz87EGR3bpOB6pzuZrM8pXev2VPs9OaNkjDfldkeCHEVc0B1QMuUb
DrU0m/928JRpdLfpxm1NLVpIl9ILkqIR40FtxOlw0jGaMirSGjoARxH706+k+HK+v4TKhnPMioKc
dmQLYCuVR6cmto6yfoWc1HmfA7AFiPOeShvfBDrFHnmu2BjPNK2gk8dLhqNs9BhkGalYnS/Rb+G+
cJO8fR3eBvoA/OsvxIcRgUTTt3vV2wPiO4YsVp434ZLAQUJaa3eWPRbbCfyFfq/ah7LK/0lo3haD
NwzuELhjTEzt0nVSARNqy2IEcBFu+pbFPB1mEWu4u3DRxhFZWiN6S24LpCNPo5ywxTha51qFhp1k
IFdjfn6MWSdbM1D4qokzex9QuvpSz6Yt6rDbEPuYW67aEhqdsRcBzqM1pI/aVb5Xhr0gboF7cD/f
e/+DTe+OsxrpKjMqT55UF3i2OW5TY3kb6NQrZh3Dc4DDWf9xWutKgrOq5ha9tf3Uh67NxkVW5hp2
AzTFjEZlKSRRW8IYR9ZLqva3UbdgvK3s7oMLNdOJeU+edM6Rni+7/3kOYLOtXuqI972frkCCMub/
OWPcb+PjZo53Nr5sLjSa1BuvDI6U6iSskE6FPQqJCEYDtQ+9GejDVElMo8U7o1lpr18wvHkoRuvb
q8c0YvPYMt5kX0NNHL6TwM9dOUL4Tj6FpkXy2F0FnqEjikaC1CMfqUOyHCczXtX+RBJ9SH1F+1Fd
f93MR39ylGyph80QBnMCdelifxnex+qRInlmSxwdutWhJj0ZnYeERNv/Xp26YDTlSxZPjUyfn0PL
XiGO/o5cXPzPypLH57jU24WIkYpFrr4ynfh6+1EY5gsJhqkHKu5LAvqsIcKmWlDpbvag4pAnTaJD
G7hK1g6rD+z/nDypB9TU3M2e2ejlURkK2Rj4QP1OzEqk2HA1x1Va2aIGToUkCr6QY1EhLN+CHhZn
yCDEIrDgfM7uyygLRsXrXZkNfR9Nj9K47uiNpmqAYgaigD2NI9V5VkAd06AyUHt34+HE99Noxc8f
ALJVt5R8iIYYLlyKhh+3uYKYRLwsQCzFJT7ifmFvShdcV6cYlTCv7PWUA6BLEBWy5XDCj9xOtIpN
dgMgbri9RYEgdnJP1YI8drqcde2vkk/oSvUXMJeBJqDq0PhOcA2l+ySNgHjwqI7OiDWREg2TV65v
4v5HVoCSy4RH/PlTfBwkuluzFTa34tIakzvexoT1RA0TX70bnBanO8k85EGY1T8Bfhbl1TKLAcB2
1plTDeKiMf6M/QZwviyOoh+uCDP0u03SVAxni1sICWuAGIlw1oAu8eZYKEe5xFna1jRIwoXW+uzf
Lip8nKF+R4yjaZ957i0PGufNM1umZuLd6Sa92zR9eab7wgHbwBxdNQLlKn5aLiQYEM3basalMna3
gKvKJIlJon0995EvpQ/s2ul9B2tlGhidiY4c5XP7eZVfA+/OYM0Q6xzg5Ggnu60UEGp9vFWmlXy2
L0YCEBu8IPvG0JFZpl0x0irxulg+Nw6QiE/RFc65QwHD0/RQvhFUgrQPgcm+sBazQ9NELXQauG3E
x5QIFU7F+7/q2ix5g/PSdAyao/43q8rB2rOHEBHDorS5kZJddzNBsxbeABnL6yZW+ykLRRiRozIG
0yDdq9nkdQgq5aj8y9HOZO64upMHXPDtcZbpfm2aFhsFeNNE4EuOXTQOzASWY8hWoD9IeGksis/t
ebCwt9tqTmUNtsoIh8sGIXWpMpT47M84TGUPCtdCsvaVDrvhaP0lTDq8VwNezMLSvO28nqKKywcn
MjBA888TQf6YzcmUexA2y6GC1W2WdV9RH9bTi7v7Hdp2StsMY32QKdQVz8gJMtVcJMNCbU779itj
1Nl/HmUfUtzu7IsF30GZos+x7aH5Odb+2UItUhwFmVkQsNh57z2yLqx6+3/ePjxXsJv/z1zF+iIt
UeinGuO1N/Pzhx4SSQ4jgRn2azgn4BQOkOsFyjP5xCr6gCc7fJvA7SkwfUpsRoLO5Bf3S1ocp8eq
Q2Y2ciW/6EKawM/y6noo/ZqXtiKI+Wab8H+/EG1LcZccuSXGNMeaC1X0+5xiwhCXVFsMxEz0tr27
0dWAjgGMvRo7LR9n19oorrcrQTqkNC2eknuYbTD/E1KQr7JL/fWse0XgKn1vuvBQCL7T7d5+bLQz
lzLJ8xSEj3S9C9OCe0JY4cz/5/JnlvG8Myi6nfWmT5uUZVi7b2cL4ucnnSQ9S1G4339A1TXPFNAy
8SZ1hMstNOWo6h5BHwMPFzlX9pznNloQ/lFee3c9lO9zlrPaI9ngR8lA0f6h2U4c0sBf47hsgRca
epoC1/jlM6QNqZJW23N+lHBUJO4wL4q6mq7m0z4wujtIKXWXijN+VZjiuU1+q6w3jZs1ClR67YqJ
X/jbBSbe+s2bx2nZPJvG7JqLi5FxE2jRrP+JPbfSK3F9JJbj7AkvJ8uuN7E0VDvA35vyi1EOIzCS
urFPWJ++vJnPF6jlYsR6DU3XcKnfi13Mt8rJ4cRmnyFMqcCmdlN6rgTqlWdFvMlSGlqhNNbymb33
TsJ3LFzrpPUyMtSXRuslVQC/t7gtNB3yZAGYK1etWSE5QhUD1hON/zfqROepM2GOZU4h8DhXIZco
ZgyjlhsEeSESDE5kZ7TaRRTTxAhEZ6ZATqaa43t6POZYLSVRGUxmNzDeUrkX3Devb0jkc5SC6Ie2
+l5HtWiXj2zg8kWYpHTIYxjDPB7C5E5kL2AfHGKaR3rU1G9AQ1g/CzlFlkBMRjIzS7u35cNO47/a
AOTQewuF8sk8tXIJwJj0YWKbwJVC82VNFegM+3VtdVDEdC9l5l4rUylfgBo5nUWEry2QRFKy3bp6
ewGo3nqVzEw5kcmOenXqz9zYnZSRKLZnBTlQH76JeNM+k6HlrzeQjiTnmgmYYYRKq5PgtEE8FZ86
+vyddMcAT1IFND2n85/nw4XLrNkj//rzi5FjHA5V4B8VHtUVywhHG0haDohnN3jrUQugOMpj1jNy
rgsJ2Q6Ye/BzZ+DofQLrRaXJkPNXKQjaM8Kc+ExNjz6pPlxZGFgrjmgb6kUeyXLlnyLvrPop9edT
A3TMwozM7RYqrmEGs/Fmnve7zJ0haZfRgKYbd96/eSe/fz0Jn8koFxXUawT//1DUu/mUVY49gXVJ
X9HccEGYUh8jXUxccwskdmrSRKus0CrvTr4CDsV/88snvlNBW2gYFYlv0AWIg8bIi87LAkGLpDUq
PLCcBr6fROfuyQ5OwPHUkLYR/epncOo/Rvfs1c7RmT953OvpQOV8tl7i7W2vgPqYTxuZLJpOkLPp
pO1aVXJhUCrUrKeQdaCs8z1m5HSMWefuWM38iDfvgf3cEIaJ7BJ/lqTB7BLzQbbpsaESY5tyQOfZ
8/nSNoNslW1/u0Lhj4mBLxgHqQKhkBEKBFK8QnnKS6XbCcUv5hIkxA9AmUmm0pOo7K12gmM/moQ/
pKeN3zb/LTeo6t5JwShuMfYdXnyfKEKrvItVwzrDLbQDxyDypNy9Qxvhku336yXHoOq1sbHe/2R7
6xPPIgwaB3VihkomdHr6SjdEjGerSGllCLmq/vdft22kPxuHfkleXRntHkTfrOz+Vn70q9pBShmN
+fTvm+5yEfihyO9tqyI7RjI0sTkJyEgWEFxKKB74pYX8HoeFFFT/U1M07sF4E4I/UvBeCkiPKiBm
YIfgvL2RZwVvRxLqrQWvwF+4g/JqcFhQIXmvs4VhOQ9Y9l38Inc/+ZklMjOqprdDGHKL2R8XPizZ
YSuukM3qCCgP/XT9BM4dHelmbqrq1rX8pNEmbscoj3N1hVQVghoaJU6RzB1w2mGNu/i70NUeLyMT
Xd/bHDU19Sl7kHktb5vqR1+Tj4X3ttBlGeTTuzXBDyYKizx9JButZgR5lKHRkc0W683LRwAGrY3w
a5eRK5E1u+qe/BjJByfsVNdFHTEiPNorcWkj3hmZVxkbZQlJWZeV7bwJ6rkGUkzqUniiix+3sOGg
xhCmWSBE6WfLduA77L8tJT/8NObL6/qRKW+/4daQZvsiFXh8F1FC/hZJw+hsC9KPrT/IN0+tDPBD
0TfMWCCIKV5ukMdBVpWmNufvcE1aG3zsj8Uqcln/tRDe1NCH8H17DtT8e5Ki5djA6eZQwt5hOss+
p7Kqm0rBWa6hW6ZezoS347opnjhZ7xAKZovSvYCIFCggpYcTjCQsqBdMeivnH8lBd50c/L87TSiH
Fpivw/g1OV0pZyOl59tKs7o4CFhkLtOUBw67zCfBlyHyqE7guiyqDZavCTkMWtyW4zL+BFLbbCqE
eOM/ZgBvg0shZFvadoVsen7G2hJRrkK9ZVk2YYDiQlXdWdrCtRA+NkL3nO8WCVdENX4qDEE/4f6h
0KTODugHsDl36OsIauJpK1+XqJ/6ITlSjfGsvn/HdSxpbtDlWqabo4yRgncdgjkfpIh0zI9s2tvT
GB+qReCoN3oIZUKX9N/TGh0iYx/iCnVNB5dO6sItqF747BNKT9PQArvoKwvDaojhK52PC8L8arfz
xEg/OLXxYrooL0XomscWV/gipyDWFljTy8tluk/lyACVHPUVmcj4x45bNnz65IrJBOmV5VyUKPaL
n4AWgdWMJM4NwQuoi7YZDgd7IwtU6XFBEK8UzDj2At+cui1/CMvTrTYHD/AaKPPPcGhZka4rJmmN
NShuSFyGdWNod2kuPWnok6DpELRRjPKO0S48c1hK6xUzfrCvQfoKPRIPXhpbBrkKiewdQeSoUg0l
wzaRIu1/JBW+sGHjNFYKsA4i8PDAy9YKUhjNvN5JBlMl53XwjThah+ddGGvVrY7JUAugetNk1oju
rOCUOqE/pjuu62jXy7cvgB21IhJKFJGIxk4Larc2l67ulFW+SAeEBWW9qzuldz1pJJ5cuWYrNxfK
XyCm28NBzd5dRX7k9FtUcUF0X3z4NqD7s8YNIfhNdAndiRiD2q2vqRhpKI8YF6p9GY4xPQtxg7XM
m6bUXt/jsJVvSr6kUx7WJ9dWvQnLf+F+uqYYVoLn3V+7MGOYDCfvyF2TT5p/GbASbsOULM3lfv/B
TdkGe1j4EfPhcX8sTrazpTs/acoYVRSG1OgmV8SK6A5xqm1yNrOS6acjTuxBw0N/ewhjb52MSZbV
HuSsGa6gyYb+nGnWOYxGS01S4Ji+0z3QY6EPPdm6Ju4eD/GIztx3ecHEzWzaSTDjct5p2WbadRxE
v1pDiiG7UP0Cn098+KS56TWliQqy96yLCgvmHFMMtnoV0IkDqExmIzHGlyf8ZBHaraLsYEiU6rt/
eGlpsr1quXxbt/gpK7fj6jva7YZOh8U51dtTYRrBTlshnAIQq+GiNQtL2D9KlYfA1o30NhM/LZ/q
PkbZ+xnCh+sSqaMbsLS9r6h1PQiwzFHDBnq1K25Aw5j/Y8Q1OamjynZQxoo/xdV9V9HxRi7CB2AF
n6f3dEVsNPo3pdwg++ybkGgEo6L5sdZ4V8H47zo5yAF7SORtwcMniM/boqPG3DweoIetFqS1T1c2
ACSzgRoOR2KVtUTQHfsw1Y6QbHWabWu8ClcI4iCJMDBWDoh6v/FQTiYlxWk/f49krqXwNws0yxPo
BwkmXI+SeZDxZnzzP9iO543AIfKTrj2ROThgUWDpfvAzS/h/RwG2QYRaqydS1mbUqhAbB0tE3agV
pqLVkZvTWfpucWcoQsyJgTsmgGGbPDWbwaBb1EyVO3iyYq6jvGkmMGx0Kj2T06FwFuWeKs2cdSp2
ZOkPlcjsCFTf69VRbUh5M440/8oDpK11E/EPAINV9eaYfP7zyu2QBlo5ZD1qmBUCFo/O1dboWo9x
uPjufCvX5tlEfGftprFDIcXU98uo8mFt7el0p6rnlmlf6iF6LIaKdCdOSqo8KeqWeQAYn3PRY2tl
+GrI+QzMWDZo/Dt9zx+ut4qyF77EWHeuX8F2dn0+2wEaT0hjSMVG4ftGaJdLkIiufQHBiP00Mcwn
nCj46m5Fb+/jQwTsU32yNqunLZS4JwFTqsd5mHRLqFLcKPKGbS6sOejt3CUChQFSPJaxyS6S14QH
SX0u5+Rl2gGnXeMuEJvTKo+Mc8cGGsc5wWzfJ0i6aFP6oPkFyq/zIrz0z3ooFpxbA59lS+hNTMfC
hlpxx0WK26oa3sXfgBd3AoeKHjfg3HxZaPybqKmmw0czTTcBfUmoyhgA+l1J9Z1XtAjj801ql3Q+
GYAAKkZslkdbU599iJetfchOD9vX+6WAZNVYwQq9uvhBwW9Sz8re4TkThI8D03Ep/0wcb3OCdb7L
iEtwIgfFNx7SOCtW4XMQTgLZ9NjArV+7EEcFwMBI7s8vKbNq170jrx6CU/MP5qDmc1td5zHYySEn
tSC31VD1PXrYxqAkGH5648v1ATFj1NGtlFXs/aetWgT+qsjD//uYQjBGCcIT7Z87QdU52HNCROT9
xfWWb8O2GN3gPa7Nzv8Klw7qu2rjIEoWGy0CujyBmMFCSB5jQ5d1/K11jr49Fhj7oEa2R7iufPCM
agHvX6qg4lHO8/K+xf6iA2CvSroqCDTmQ3P9Xv9UOP5YUq+KrPfKz1SaisTvu9LQtvegn2M4dcHP
4y0Pd1uo/ZIwZi2Sm/VE8DOvwf2sew6cZyZcIF8OOM7Oeg8OR+OhZUrJJTXEq89Oh0Xl3PpGfntJ
ETQwMgfKlTKpTEvQbquUVrr1VHEkBGvEmYzSvsSI6N/z4y71YF6Mou7CSIrxpmvGXpE5mpTH55l9
w6fBfTvudFcZsm2zXUfPmqXOLEATbzQcrzon9imu71t7aKX019rHHw0plczW/tBJrnMnupCVkTwa
0+UWRDpgTHP6mTqrYNFocFA2LVsOEhux1wbkgIvvXr9Grpc8X8aJ4IDRHYYjE3pEAYNUF3W3h7kW
lkgo0Eg3y1j1AWL/U4ihpZVzkwiA9XEeovYuDY3g4/oi+03GWQdfw0GP6hA6GESkf18GjF7BeSu1
+cJlXOL5qlhTathkD81xIuQCzuY0OMzOHWUsMF7Hb3u1vNIrTqPD7OqszPXxKN5Z4WMw1qxvYd1t
u2edezh6c9QDOGlLgM9wW76eKka5QQtw3tXGBrn+5XNl3+mXjDCmlc8jmoPVFLGwVOTo/XAHyhvB
r53Wt/kKx2kocA+lh5W4AY8exB+zDH0WmeLd9ijF5Mrbo/CXihNUwk/klSOqPt8AOMoK3nDbf9lp
ERU2eu/3s05shQr/YGqsobyfUGVZV36u+NbjbMdj03Xhy9iYQcl7QkaJvGdoHXvZB+xWKc3RQ4lI
ujmcgjH6UDytMJ97bCsX9XP/OqxJgbtn7JBYFTKVMYbNoD4ePFk9tAgfQfjlbY73vX8DICjV1grp
Zc44V0ubrIOobYCbes8D/Y9rFbD0nDLijWuJ16K6zkBMz/JvqAiqkNbGrXqXppnC7Zn94jcKcJ68
W1dzj6K9IKc+v2VYxuS8h5iz4vm2+GbRQK1WHhlwwQFrpwYUmOLkV+NriCZIgZxFKOw4EI+SuQsQ
NENbOzhJdHyzJP8xU9xcVaqgq5AALBRB2qzSsdyCLOPBkuD2wqBTBd+jMbk4RPGghcK4+ToJxImJ
vFQqER0Qe5knBRKnJuvN29FcJpKho2oS/WGx3ys/zojwhi4WUFgf9y6DyFvR2VSI+AjcjjiXJwyj
MlD5wz8PCCp6sSi6GeIpF2WhkAm17ssTNgcW9YEX8xFRzqDLn5qRFPyERRTjuc8i3sNNh38O4Zkh
WaE5l0QEcRuJ4oSpoKegdc//O6DsyISsKCkigvwH+zswbZx7goWpHOtwcm58OAn3AvjWb5ZD9ibN
3vSQya6FgEuZC6OcYWF1cutivcjv1POANgrqnRSMDQPmOMg/zgh7jsPSQ+E18VndQ783AWMyHkUc
bUSiRKHMAgIE2PhFHKGVDxBZ5Bz3lhzbt0NcjXW0W4DlSXbxewXD77464GbwWQ3rltR/e6m9Mk98
ksBObQRZdx8HY9dSSHJvKw7fBdJkaGPJ3nOiZGKkOkU2gdrRiwIAZe2a5AuGM/Q6/ZY83IiX4zNB
+4TjLQyAzUeM0YospSQvBkXSsrnGR31raTSgF5RTvtg4mHDRgi8qMgFSvTr0qadDb+Q+4o8ZaQyg
p+7fNTH7IYyD7P2mHd5l2sywKDflrJLFdDU2cfKGOzUbgoj23AjbX6MymeH0zt5Mb3KBNc817POs
tiwkrTDqyFs4dyYnT3QeOhdp6M8sSxvhvtTaeHccVvyJBtd33q5/IZ7GGP0wTeMa+HJZjcRUCQOY
WN/jhHRxX1SbQDkvggVEEK/fQpmej0RCnGhHaPOSZ09d0ruvZ9KBl6Em5sUbp+nt4tpbHdhm2fZA
11/XAMFqUlt2bvcSoMHzzENFb+jT4cPigGyTjKN+K6rgt/N5KxExRjBXiugzKbJgFoeKwLZSpkGk
AYVRDP77ATjBADv9dv13q9aK5LXUGGhC7I3raK4toYBreeDAXFArh/m4pySQPs6oafC8f7NyBA5e
5sONP4zwYQZrgQDo5KanX6VTg3S4WAc2aoiQWSoB82F1LqS5gsKhfmgfB9PYHR8a2rH+DeO613YM
cIitTiexyNrbpYtOhr5lxZ//d/FSRWa9jsHOShLWjKS8LXnvyG/5cQoH/pvnkcqDJWz6rDEujmqr
aY833uNyTbW87F9elGK/Ys1u8KGjSx9z3bn8UUqVDondvZfm4PJZiiSZIMFUnYGQcb9EmZbu6zRI
HH3W+v107LCPJIf605JXtiLR/sRGL0hDQUkiqYG8ZnD5YBUawQesDS5A7sFV7vFSTrak1QB1O8/V
FSASU3nTiM87p+gQ29T59CP80dS6QK00jLMqG7jD+3HVavzv2cSyMv/QkGeR4NU7+fK6ZmaQBJiq
gKmSqpn3fZaflunRAwpc8l754uhe1VQfo3nupAvBs8590lN/eGcsshnMAvxRomyc7mjkvzmHsdFy
r7g+IB7Wyz453oWVf24CCetrNMZgKfl22kU+Vfrc/ldtJtKmD3tmfaMxSK4VKZ3CHSf2+gEzvo+n
nwGqwSZyeSaa0JnO+VDCfMmNLUlaz2igVIYv2kb3osLhDedg0PdifeQryh/RVkaY+0IY+3uwk+i3
bBswbOCESj4ZtvKgRuzb7IHpe6e1xyG3Y8xowIMG04oWc8JKj4eo1cEtinEIlFtY5YO7BeXn4Va0
8jIMt3KKMtk2agsYe8wo4FZfGrjrxFGPvM77TsAYNEhSAvh0y2N5G8ci2rSV/WH/buR2YHenHDTw
oHKb5ZF6V7zwcM4KnWiqXSWr2nJbyNhv2DP0SD6w8cwGclWF17kyY3KiWdEa7nnKScX+8Jb49s/8
4524W0mLb0WXmkXOpQSd8Zu97p1S7df8CCeZMR3M4bj9Zu3kPbdiJ/9QAFQtuRdCd2f7LlSqDf6a
w6FbMjWmcqj9k0WU51ljo7q7HJy2j38vQd35Aq7N2m4wseusYwe1eWGzG3VPzHq5r9aFQ+c8BEOi
TGxQ4Gp8aLXqKkC4dRHUceIG0jzc2HsPtrDCH4hPFblTcD4SzU/GUQgUVvWJaNgXssnFUwFICu4h
KnjTPvwypOOl0KzpyFAn+qBqwfMxaS/xZ3pk93pez+2Eeq5nmHXOCo1QM1s4BThHKciuCYOnTgwy
KCgZznhSzf1w79rI1ZgEU8wOUG/FLHxWlQYOaLwjAtConvAx60MvvlneEZ0ut9XF1ea88bXkztR4
UXMuEw8biEw2m5qsHANzz+yRqXYeCmTwAgpMsei8iIsuQUWtgwtMT30cOFHb6gGgnpx+ZW+Eye2C
pVz8yNeUfFhhMi19WJo+RD8CcmsKXaVjjYWLDuFvPFjnrUtX30Ch7t3a5dBS/a30oC8TFn83ClLh
3D57p5TcnbGU78JqSaxkfinO+nL5b7GbHgfq2CHJixgopfTaTF+NGfUaUyRkl98FPmSu3hRqchkd
ccLyjA2UaoFLywxquvo0c6xbKf8d9Qx6e8gHQAQ9sZajT3y79kcJ6D7Njw5rlmReCamKiHembNH4
LlYheDTMLHUkPzf0moRSKo8fV04RimdgTTBC9BfGJhkP0tHwRs4jNqb5joTLV80cGGGFw5xvbYt9
BFZowSG4pjGaJMdPmHKswpX1zQ4nwe/8qT8/LduAW4Cew7uM7/Syc/QKSXbsCGfCpGCQsIFiktSB
BA9S1IxuscvkdmiKqfBk0vGcz2pQ92kDg4zxipj+2qPpgo8PJvOMVghvQrCEDXOTkm2VCv7Jr15J
Le4Dstei1LloGcw+qqV7lx2ueXXWOhoN9z7dr5ErzvCzNCfS3eEeD0BJ7xG+J7ID9qBkBnBBdY83
EsbJ8SswqNr7fNownEPXD9zWVs5qFQudKC9SPMCej+Am/LS2cbBABN/tbU59ms21iEeRYXbtGdye
z8qPasbCJNwxS6TZYrzbRroQKJ6bx5WoZSWLxbiZpU63u5SnVyi7G0+9WBlmINCVEih3mb7jiXU+
Z5NRqwLUJBPYxqOyef8IbhpOP3pY5xrUG/nyfVssxPmit2E5+S+n/avV5fOnIqN1YjNj/nxmoz3Q
ZUxlWrqftAcxigmdloN2uaVBRTVqm1DoTJSpqt2zHiMDDV2jeYeLPg/MW4SEZaEs4jS6kru9OjzP
FBHpwIFe82nbaXxrrFUarPqI7Ifopt6z+LD4hkbusoGEkENP0VnImno6fLOIz+7wVKdpwtWQD15h
mxz3u8VyPYeBN+pHWjSIdV/b4eqB387szKAW3DG3j4EM3dIqDmzOdvd3g8mUEhULM4s8XmatwoLT
JdWjMvdUdbQg7caVNMIi9gQCuXbUkF55s3C/ewphUPGOBjVqj3jFQrxl2hf/s6CnGdmVzlOHpmNQ
9+NlUWAnZQIewwlZiZ1UQcJSgGqTDOdw6iwtAp9ejxb5/1AJHEv/cvAM6dlFue0jFSafdLOGSIG3
Ev+XH/mwOCWTkVSW7TtK8lcnp+9hC7u2kSEhAXe+vSmZmbeoADXxXImvlPzxo6n/ob+xjca1vPmE
WvDFPZ5pxcffnliYOB2jNtBRYk/XwB4l1ZhquHBZI4DWgdyFwGStypix30UPz/ZkmfFKj5EFnFFu
UboujaQSMSv7YooaG+VW3WWWBit8BgK1jOcArQH3+oHtMF8GCSRW2NUOLY3SESPMJz5VMap8DY0d
XjjYezhe0laAim5wjaQLdOcajlOREvn6eiqI5iburJs2qiOrxww0a9EJVckpMAMzwOOipt2+7maz
uuJo5i0vhCcTSTQ5QV2AdEDMxFQQwut1xYQ9C+JF6mZ7z/aLVm4P2h9QU8Q0KylIQXMtSIw6Phx8
6kCb2DR+3neh87WZfyZd4neCQZ4DOUrwODrRD2eMnpoF5blgzHJJQa/1lvEBSNakmIlIryWU5va/
HDMxZ5oUgXlu0Hf7TBb4OqwAIfoTasj0/u4uD8cM+g8xv0OxG9wwX3235tOt5wxDO0OUlV3QLqgX
quU2XukKCxebKHxtvVJoLxeNez8OAkZWlEeUABGJJoo6j8d7vnC52ma0KPwX36kuQ0DRjZazPQvj
ticABMPOiYJkSP+0w/eqCHxaYF9kVpH+1fuyHCaZSb2+lHysMdJKayrJjELULhYFDjzIO2yijpkP
MHSOseMKTirZNHQDRfpQ1HKKwWJ/tmIMurJrjQS+j9yhwXXhy53z8aq5QK6vbRUFdtLjGeBLNume
/wSsFkKrxCe/7hpVL/nFMkqmXtqxKMSOo/OY2oRqjJ6qCU1mex5Om/8jYBJTSdjB7LLScdYCC94H
KYgQRSsblRU0lbrH70JZV42avHFPAKQrPaQz9mK+pCCwxvmqaN2MLh6spLKBIQwXoSYlkYAmYp+O
AF+bH7Ylt6+XkELCMlXpSy8aJewdIZ1nmdhA+bwFWCqb6DtqUVMWB+pzDFFz/o1TIW/mgUSvWKpX
BTVXhVyRCYjN6mrtjZLq1KqfP82iWpGHWJH4cpsmVpBhph9r7w/Qn8+/tZVlXfaJyR2EUst229LY
NiITjyLBHP/b5QiyJ40AeJ1+2RHFGYoajbpyAuLDf+aqKh799B4DaIWSs+9ZsEiZxyHeM/AQfwCd
8I7HhK0fonxofTIBYynjSxJKpSsrOi7hDpgxLIvmQm/BXLaHo+TXjCsUwI82SpEeOSNbbSKTLA1w
u2M6kJmbMNIJ0Sk5sbSpaMbJJvmd8TBsw57mq4HE0eoxWQW2UkgIvjWn54GxilacAxcnlqXJCKZU
dmK4krcBGkXSWR/D5Jm/yM1EddnuPHwOt8h/EMbt0mpGWw3iWFb9XmeRmxtXEaJtb1kXcW6BN4lb
/yC2nAOLCrYadoclerIgkNgqmmJ95qeBRLOm65256rpXRAJVaHrUb3IdNNMRJPzjH0FI8lybyfvY
yX/GkUTdrRe3wnzPgj8dn4Q0bMZwcL3ucvB6n9fcnJvE8as5PRqeuG2FzbGGXkD1G1pyca3jtFmw
FXukFFGN/iC/pEuUlG0lXE3DlLMN2YRkUEGxVaDj91cQRrhM0moKZ8u31msTa7nmIvPi6aZ9Q9rx
w6L/aHjVt58pX2/CmPSUA4TALsKYKOkpt3uhO7qQMuXqMM3HUZDoXxFmqlbwUCFFx8xRN294doXb
DIvtG3d/l4HkIVBB+FXBlGoVH5H1qbok61SJ+omlH1O4u1AjWzLt/xd+QfqcYmFZHEMrJYunE/tc
EzjmQ6C+LQyHsfevCqnn/FiUrNle1FR1CMFSaqrHPSOgno5K75vSClMSXaNn1smDwokoGUzXpW7k
tBZkF1UwcL72jJ4JF33FTGaqc+UIF35kN/+gza8vKE6YdV7Gl5RpdSpUgxq51ltTK4RmcCCWg5q5
SsYJeVOa6P9AiWsjUOil5lvvCX8/CpLlHftZCdx5NpX1xEqdDCND9g91HhtWEdqhP2kIqpnxp7vY
yBV1iruloSPkXLxKjf1iXYbz4F6Xt9OTUbJRG9yvFyr6ESze/chvDC7EOL1eIKTEIU/EQJsw0jgZ
aGWy+hJo+uveruVb8dqVA6ww6RldEFpVm8QC248cFA0J23RGQMJ292e2NQ0N2maHGmttNke2aJS3
d5Q7rPOn3zV09ifIFLWsItlpPlYMxnNlJ5SeuVoaZ9ZOAZgeMknCIC0UO9FgaikXjd6vWtNnaFOE
7baJHOgmjPAjMgE8p0S69xJIeRYBSgaOwV8pW39whpQ/kHZl/lvUUuF6gXIZuCEVLnvKtE+Eros8
NAP91jLo0cwExtYGE7T0kzB1XPDvZDkzstbzmj7/io5N4OgKixUGBSuguc7f1ErdoapM15GXM0cD
KXkHJDRg1n9cir3Ngp/BTAHO4BWhwuNsprQeZNWOB26/u9VXPLEiC+01lMXtlCkW6XxEaXbO387l
x8knw0pxH4kFiH8f40Euz5+QGhx8F3vIx0vXNxJgBuvB4c24rnjHjFW795a2TTsZhc9NuLXV5rWg
UfQ9pK3/i/0/FUIUc+N64RBgNzDhhGhWKCV5OGZfISjGkhBdvATrz/Nvld8M0bNIQIUCDwuNyMGK
qMIaXoOOqk+4huqd7UG8X+bLyruG5yzvvcCFZs/gs3LbviZb4XSn9GGdSFP94pyjHsjaL6oligHp
dDV+Iiw33WN4jvOQqFaTNW5n98YG6kSzmD7mpW5JekPP4yR/vMEe96nMsZVSjmj8hQOMrq/KVdh3
0UH2WjlOnTlKNsoGYBkDpL+K5ZHd/lZBnoIEbQ/CThEJ8XcD5VeWpMa9HRCSJSAaPjcPg1GnchAY
jPAj61Of5/3VyLTTaWNPHY4+lcZdTmITUgj3B4MsWWaPpnLgosc8F5wru5utFYP11c2QTHLDGoH6
C20EHhqnX3boqgPmZoUEjX4WBa/n8jc9zMEIlxdrREwgVnlIl1sjC4lLptbwjwjxfGYU8zwizNvA
RMEReUIGryblERp8kB85VK3Q8ICEsxsHBdROUDCY8B+KOjeioZxFw4MyIO4djj2POqLjLy2+vFhs
EhbZRX7vUh42+rnq09653X7DKLWxt6o17q2c0Kvx2Eq/PK1cZUKNyn2X/G7jac7lho/E1ZhvvCBg
GxrLVq8Ns8bHRmgZGUO92dLvE2Ja647DzGSR5YGQEQES75vlJCaE5fDTvf4KQcJhotbGz1Ly24KD
uphgJEooOdKjhFCbf9QdeMyfkowZoCcKXjqaCwzLhktGIlqOePnflhC+gnGit7FTGam4kqRMsPOz
5u0btkyBChPGgYGfr+R4wZgShvjaNEpNER1veI+LZkVDZLr2DM3sH6Han3PyIZlcFKNMa2up9aWs
O/dGcRpGx9BH/jLcnGvYHeSZjz98QlPst/7Q1H9UGRSkdSwv/7P9QWVdIcNoiiMqTzuHJ61AEq27
+wdXEGs3YKkpq8p2l1CqGWGZ5GsYUzvkUDoSZm1H60XQAojeo9VM9dRA+KOfXchvh3CRpAgMmrFJ
djyyw17127lViW1sohdBUtcwUyTpvg57BgcnTor+bLpRxctoWn8kTVMEam90bJz4l3qoyhqwrT2i
nm3A/IaP6y3+ztJV49pH24ltiomebdcOoJ2ZgGnqt6GPnGiMDGWQDDC+X8UEAVeXj6pD1++VZnUQ
AXUcVqRezx7lYi4tpMj+BfxZbrH65gsDE+ghjOXiJSXcpwj2qM+MSaiNlAgMykQTFkz2V3PHaO5f
adHKxnzL5hGO1j69PI5/2KABO9ljh24rPRweuO89H5C0i1+sy7Qu7gE+o0nikMLu9wFbM/Yv2kjn
rYWDnduQfngeEBSVnH4qADtnd0I7nqAenWlElbUOcvkRiHNyNiZ10LFYl7QnWZSOi4B0vZRpVY3N
hAb/zLlw1GfZXPMfixumjkPPGpWdBj70GG9qr2cdnfmBC6H4Lm/cnC3k69O2swibRZ2rkFMuNQR3
bjymSpAV6GtZMaVcWrLqJGIL8QZaRdCYwWOVqj+PC5o+Bm9kACw4Ou4TT+rgBJv08o6hSB5ikbmO
qzKgIdB1VAKyFIOBDohrXtAJtmVlSMJfGFqvuSiZ0+MgSOag12TvPM7gr66PfYV8JkNAp7uOWyTz
twEzDJORQRn4DyTNnGjBioAwPLyxlXeLEFX4+9l7si762QFhu72aQdOsqHshMr7rQ82UoqBijg34
2IfpiW/W3Na17GNfPmQ8QRp6o2RLUYML44pV2ncSDLEDPbn8wFYWGwrqA4PUPjiD11gDwR7B5Wd2
AdQ7d+PZl9pq0VqmC3MqvX2omA/R+qneP2ykkEoWGv/eQPa0iH0wq1OdUxrMChhlt3Yi1idX+3p4
/i3/S4ifJLBb3oy24jLzkCaeQ2aBLp3bSpW7OAPAJpMaWkV8TEeVEarPDCP2tgEx3Q6gkQ1s7zI2
biCcMCfMJpWh4Z7aIUcJOz73pmQJBGFCKSgvc6yn7Tkw2ly8wct//mmfbcrHW9GGachLDlA+rvk5
by86GFzUm0A5HuGaDofu+9q+/ls0hIy16K2TWxSgkmnixKmYp7ixvUURheOJy/r+7+tBcCJzvv9k
b8mYv30lKTsKlr/KLLfUVQPRKwJ1maEfOcBu+BkO/e2CIaKYP9h5SV7ZWJEqKycqCADHbC4WdK9G
Iwng9xHvNeddZHmSnTpXyVbNT/UQU3igDzMQRTXy0NoWZ5tOz6y9e/Dk9vsvqpdEP7obmqF2k0mR
TwRrzsU40TXWrrjAlc14EF5WAijoXYDzQiKq8wT+nhhLL7V+qbLmANL3PRIc9KtQscw30zDqsTCp
/Y/nevlSO/GdmzsFGK7+WX+ZLKRQdigHRK7j2HsjeDMI0z9WekXPAlCBSNuJp8UvwnEBdFZfnNTT
+2nTkfD0MklhPvzf05S1g4jteItkiNhFpq3JjN1eW8awSh+NsiFq3fq7FT1fCQNO66N94MmOMoEP
0vfKIspid5uvL9m962MzYgK8U8Jqz4HkyRPZlSvLn7zkgP56noCiC5Ff9Rrm0gGDu5GkZHb9MESP
a2j92YAlOlpICpCAoaEhqtaH9aThcc5WXhnR7u6YPPcu2ztIOL5XF10Ka6bbIjNMfLT7UokwckI2
TdcRtWNYuJdb23qmvYGjbpFEQAce/ctIK5R1b6+P06nGYu+N6DioFYK3Mlkll+QtpD5soYuwOeEU
gKVfzhcR0iIbUzlJKHKd1gYtLNdsZLjRv+btSFWfGEDri6AHYxokUO8vd5ogrgWMZGB1oWEWHgBE
j+112aJvS7eFQ7g266fw1luwIa/9VxZvBdNCX9nu2VlSFxZeQfN+Wv8JQnjm9ezXGyvbG1pooZSe
rpsPe+3CKgG+/5Y0P1uctQ+xbYxNyuKWHxaqKBasRQGfzfmJvfS13KGnMKs2WcnWzyv2Ke8kcSy1
pjnHqG/9NEIRckrMpDlwI1wkOrIoR9yRqmWF+2uaKq+vLu1sFXzO2cvtIBYgirmQB8IU+Yw3NKmo
KUdguOH9/2h7vB9bBvOI16yXCdmCo7V9G3SxoMhqhtNs3gWMtgliebmwoDa7rWj57lN1AdmkD1XS
ry3GV34rPe+MegnPDfcAGTzeRSiuEH801gPxc1oph0aC0etQRKesLmtwbP2k0oFmKqPbzq26Efk+
uHreB+BNPVQy6aasz6Px5lLvhck7JRRnw0HzlAa4NACH7o+WgWu5IoAk2lRK2Rb4Th0Tf2DjJavG
adsVEUWitQF/D3QZdIGhwbNisVg9Dn+BJgEHJFxmWRAOgwEml2tBM/zdHnuhsdqNlRwVXzB9N0/y
m+BXPRGrhlSbc9CGSSulRlXSF8+Zj5ATwSNsf+RTKm92g927DoxWJY18lcUT3aO6GKDkbkzV1KaS
mTarcvaEOPvmMSimYb88rX4t2Jga4xEb+qNiB4qdnuYCtgzjAuE/1oAV94ejEOnjcEPzSdN/t/Rn
xysqXcF81FcjuTG0BIOtXzGozqqLe9DpZEdNrlVLgCwbCTDG41R8MVPXuzsUXZI0N0bo+OUeyKIP
hyZ650jJHoz7/CkXPit0ckcrm5Iu/j8+/XkzeO1wwf7iJV8h0jHZD/L3pHrMx4OLShEeB1wpyzUT
vNSO8StJ3ynjGO//9oML07VzJefqUXrOhBjLdT1IlfBR3k0wSGSskAaBA5W7Gbylv05hqp8+t5iz
8RnborXArSrPbKMpRobw+rhUJvBG+JOE9Jz8JuJCSMBrmVdgCIx3N6u4wN6wmaaS5zg1tpoJnHUX
mEKZMcH695Lv6mO3FGyeXQgDfa8gi6bjs6zXuh5lwdA6F6ndLx7pw7ujsJu3QhR/0o5t6i1GsDsV
xK1IEpUydmxWqp0ZFkQwVD2KjYvj/CrdlPP6VrIIieHvJ4FFq4/EwfcV2MLVBi9TMg4br3c2hyG/
YWjX6bL2fWHdY/BKjboEHYKcp8ClnBp5x4InMFvA/z7lIGPH0VvRKJV0hebvTR/WOGO79b60kOhL
/7Cq9WHX8dvqfeJHpuwOHWzFK2n7MjScxMsFGVhg5FsZnRbcPDUKUnuImtfxBeZ9SJrDUfjMQFOq
qL1R66FkZIpiJ5JUR2M2Yg8PN9ijCwvNNZ5Badl3lBf9TD6BV0n1zHkudTb1mKc2mYMWi76yZ1ov
aL7JOd8Kpts4sE/3b5RAS+cE7fJh4qA4j916bzBGA/aLNulW8amo3hHiR3drq1T0VKwpnh8canVr
yaf+0TzntC2Y/XKmtD97XA2xHltSlJ1GeUOOh0X1PlW6mARM+YsVEoD8pZLSbTbFAn5zpCSt/iCH
IcbeYBRiwTZww/A6TvOtBpdL0zt9cc5sdZbeGloD62snGohmtbaIvX6ofB2x4+Caf2myZGroTU0F
bYnXqddofYSIrf0rHtOQxkC947ngWcJjNgH/Sv8G7JxCcLG57lde3HZIwQBhNWB0ZPLE9+SdInuO
iafbJGf0sZ6IgMUURC5Xk4SqMKV2zPdlPEVcFNZWlNnBhNVoGiE2PsO0j9ZbtNfh3utMW6XGXedT
+eun3E4q15RpJ6JGO/Y18JqDRCczWCorakk7CybrEnsA2T+1zr21lG8jSZsZdwrm5evUaSP3sMpz
g+ertgeAWCnwwg+DnUcPi2pm+p3JgpNGa6Jd8GQVgWCRwO9xZ7a+MrhmrDs+d4E0HzOhDPBew1NS
Xw4rVz1s5jrmQG+bAy1KzBn23OPebVdRZgU2sSk2+ak+QMUc3wys+YFBPVqi++gTCNeoV4xfn4w8
/qUgsZ+KNDG04mlXu9KMxB2ETwlp2HGtBaPyIa/tcDhDkAPnVeHgF31nKmKSufE3PnJxA2VKne2w
8VkAMGs+Lul91aetcX86YWj0S+67lRTPcYNwQzdrx8jyRJSwRA2o1LL901f+iXSUxnshZlXPGwCM
olOEIk+sGmQ91TPfnketo2SSjKXQQPmyF+KYPCjxzKFhT7CGQ6wr2NkahRNLnEoUhsWuX+jnHfKP
yvR8XiBrR8fcWKQ9n4DRsYY93tdAzJrh5YdH1ZcFKx2JYbHHIEw25GPKqo6mRbMCEtEgvz4p+fb+
F2tvSR0IPQq8NmwaSVlJYmPCD4UZFX8u7R2vL5vAl4acrc8ZAjNnj4Fl4weFpl8TP4wlAzkjiiAN
NWUskbsprGaxLrUT18zHQR26ecnSL0TFeMMJzdyOnomk3TeLW5vAJjM0hsS44aek5Lb3hTJKsoJe
rDlZGO/TdaTOLbNmGAfczNCOCjS7n9w9TNfLj7SZwWtBb90BobiR5YlpE2tKVCga8R7l5IAV4pE1
VqMo0ppPfLU56Qhd6yiCSflzveUZ1J9d+inC47vEB9Q6hOEtm6bOSuJoOyGZNBMK8tlF2G12FOBw
JZr1ouUahnFdaSGy1Oi97xzH8nZzb9qAzRsbmJNn8n7LpLzkK/PxvzHzfHm7y8d0KXdliZ7aBsMW
DA7xg11fT9QJ5Ilkt0EiSR/G3vj2LGdVQENOnfPfuov4RLR16BYG+TUwcNxBiVfegyuGH1f/HQFk
RgQSOtGrEb6pfURYTH21XhUNFJB4dqR7TVKK7oIxAhPlGuo3opvOvOMGa/mOZh0Fz14nh7ocOzpE
RHov2Xy/+IfZNiK+KOBP6G08hlvYkN2tdBP/+hoZcLGiLPA9OjbTqP1Igz+MCEMSJle/WtbgSjrx
88xJbSM2ox+JW3ppBKIQWlCtxdY8BLKGaCOsXbUROSr5YE5SHmq5keA9oomdK+C22oKMwNJ0f1Uj
UUgq7iKtNJ1lnRHYol6gaxJhgW7qGAlUUlZ6zxMcWW40sXpFk+kW+rrkyOA/N2GumWM5gzjk0I2F
XwoRJHWcd6qAeT562UTZe9/c4pcym/8BICng32QcTyja74VQF16lEPi2CubQttLTre21/tWvNbzi
Iu6nuKbBmGeOlPBI5vpHPXDGcVOFovbOYkTO53UV8ijbOavqHDJL9PU+LLtg8gaudIHxgM5s8+X7
r5C1PQHDUWAvJ2LUvrAqpAoQjHvmVO0UqVHsqmxbjCbqKseN/PeJ2uprdyEE3QXRcX3giHdBAxHx
+L2cVkaBMdbSPNYy5EVXtoWVj3G9nB9QqjMSuvwvCRLKk6Rc16rFEeeSybchlAHnyg6tjXw5u0rw
OOmxjwB6HiQjNmL8tCohe2M8ppvhHFWYGvZV32EO6ILEZIO1xJqZN4I5vKBVeiU8hVwVAhQguNiH
1jzKM04rTenGj2XvheU2uRQ9r4TDIaHvDKlrKVZgm9Zr05w3hViAsMux40He6UW/Yq1ZWQ38nFVd
2KtPA8Zqr4JY1JlxALV4SgIAglskXVQS2VA5O83OABFaTcnq8irzXyWZhfUsbeBvCsHxaiPyogaF
dScnAUcvm9wd2lavEyvYU7FFggL4zDvtrI5KqPZxGGZkrtgq2QvLZULRoCo6O7l+WklWCgFIfylO
NqCFRu0yvOcaD1Qfa8/+M0In2BqCXedBf2hCXrWhYuJH5BG/clqX11kdUxgoW0YeJwYKLiCi+/Eo
8d+1E5j8wN6UrQ9N7921qlzkaj72+i8ZpJsHypQV28twKGuFbKhKFg2AJDL+0CoHZI3GTSbEfKMs
ERKmpdaseOLmLYXYc4D788kLx0J/hg0Feqkc5lOzH2959L2Dc1Ee0nYVOITLdP0ZaDEwpw8gQX/B
z4FXWOYieKiM5gctPJT24wy3uNLDKFlONwAXmviPuDZGmKug5VB7wgQNqEuDs5CTzat8ycHYclzX
zW/rqKZ+ZjOYYi40jc6OB4lGI/xIV6yLnwTw5GgBaw4LuXxdpAGm0lYxDVKDu0giIpf2k8v7w5xe
Bpz6lO7rN2fWc5GGGZ2Tp/zrm6BcX1Cxbw6IdSwT/Qv7qF6txaJhdCCQsxL5VD3eupsz5AiXqdpv
yOOJI9Tsb7f0HQDdcHJxlOkh2yTyMZsIJZUt05jvZ0qkxzUGyJgDpZagRDj+PZsXXPuMWq9SULHc
xRVOjIEucGvPGjREsmEU/EVVDF1yAkQfqZpTUa3R3lYLbVRQFj7/HPZTwOybqI94ee7vbue8TJK0
v83bPbfN/pEs1fi253XWQfPeAPH4wYdN5t50CR4Q+sY5NRL2H4d2U2MFW90OPMvEOWk4W4bxhgWb
yExdFvxuX2OJCTImAhWR4TxpBrQsXtg3FJwYxcjB0knI2HRp4mYAGR3Uoaz0VG/WAYStgHyvbNaw
LId17E1ucj6W2VrxTNNHLt0uyng2rxgee0pbGATv/hyOM6rEtGEt6Ib59pA1CUBFsvenUfIP47hL
JrPkvlRlIdXXP7kvy8GtAUE1RyqDCWfD3FSjuy26ZGihooiuYygPFXw58xRMUah+PSDiORAWGJWD
sLW3/Iyd6kd0T3pLyagYYE4EGRM9obpJKkmWMcuBYC/dyvWPyLfb6IIb7VMmZXeKMQtXVJY85Kfb
DB1MHQL2ykwFkp02iC9pngt2diOMHAK0HjAo9WAxdfxqhb6r5PjEQcrp0TXUDMk51FEUfqiXfZdU
wjQRUp4oEyPgU8tEZP6Pfujcs2q13Dih3ZkCNENTmpqrepzozoXXX5pTUK1F0FfxZY07Nqi10Rl3
k856j/clW6JJxFsGpdsihpbGQCQ9VHv5cT4M0QY83mn7WWBI5EC+5nvxQNJrkrLnNZGWvO6foRA/
8WrFdIKdJ5G420e3exwqpK5MOX43bHGvZUWDBY4J29KcMcd1B9dh2EtAUUWYfVLzVF7HJaMPCBIP
j7MzRrgiSg72qSabcNlr5RSwc0x/pC+DYli3pAZVAIYWZCgV+DZ5mn9d/bqqkumjIaH/iAhIUha7
DK8sfWM65U2DeDkdE+TfA3ot1BOvQXBrEeH4SlzHMvu7EYW/p5p9j3lC1yVC6svDZmXu5y91GmRX
XyGj23YCAWMionfPja3oflrpmNMuRDkCfCOGgy2wDETPkX8E/SVOZLeWkA9MvyaWIffCbToCzdIw
6XLHJWOicVOpfrG9qyc8b8jbGc0vJDrfr/MHk5/3oBrYNU79UAZfEfL8cv1dt4XucmQfHxADZ0g3
cziS4JjQiNNicVIB1/nzRDr9Q+I2Kun9A3DT8zfZeKSBbygLU/p96yiLSpc/dJiFXy/EVZeonJNN
yES+i8jlMxBkAcw4RE8HkT2DK4o81OnXEsxRh9nBHvGiJvxFWNwdZgT5aEt/EYafw7gZXKKBrgUo
ii3NK8iIuwa3H9DcYz4El+OwW27T/MA+u6nG1l8UfRcl4Hww0uPyvSrM2d3HsHCbr8eua2qQkWFD
tyMmt11QGs2ezEmLq26cb6SA7F2bWJfSfqCTjMG8i9j+70OPUtVENOZNtep0xqNpfnbZYSqRRIty
FWp2f+GuWmtZTu0XfiWJT/Zj1drDPibe8HiTq+1SwA+1IW5zw1YJu2j3wrf4BjgvVz1TTHTo1KPq
EHWJiqnxDG9Vt810869dQcoIh3NgFjkSK7oep+pvMpRBtsF9vVDN4hr7WJNLw82MTJ+sQZEr9Bjk
km73obixJPA/oZ3t8c3mDQN8Asbv7/px9dOgnH7t5sbX3T0Dwtyy9C0Ko2gjusp6fECYvh3jRXZi
peErmUghH6DaVrHM15BSgHJPlxZCzHcgEMtOl+SSUfZnsSAbWWliZ7csLi7K0ij+m7UYc934yMk0
i4vOyE2EjR49fTPuQ9YeCkTxi0zWrzzC7apAQfIxNox7ztiKhIHO5DI8RcOynxo9tlgsKLfXLT6L
jmi651Q6NmlPY2d5OmVIvbmRjDQ9MlGNHkSKEK1r1cZ9gA5ERihln6Gzy1CfHLLtH5QEKG9hosTC
V4docoCzs/TG/v2EsUemuxM5D1MrJ+bM4Njg71oNjP3mvsn+zG1cioB2126wmhiZLONVzm+X6xBa
ZiHxXOdo85JrnA2zdQazjic9784NrM4MpiMdBPxj5S6H7u9FkGLcYsHVJCmX+VNuvkN0I/oRXOJd
TdZrgMCCSRZjMJ6/MWRUB8ArCMTVURUPOpfGI6lrtS/628XGbLG628VFtEY/jYYxOLf95/kXdnVM
fKH11UrTzSas1hxTEECS9NgD6iHfarvv0rja2xgrIjQCW8ZCBy/kv6IvUvwjCFMQHEc+Iz5AdH0+
lTDg3QmiZQZ+DFOiBRZ01j7o/0u9fb/vKarw04w9qDs4RFvBcfyis4Wq5f8tI8PeuLXRP4Joz+Nv
CbJa3f0t3Mfw3icMgHlxmqnHIjHDf8Q+uYaCrlSBxX8KzLy3NgwXX0JhlVRY8Ut3YY5VGmx1eewi
yGHPDb8yKzTqFL6HKMUdlxRm9e6DchQAmBBK7Y3W8vCg/gbpPfiUOD7K8t6PvGxLGdBYSsCx8clb
C2+QuDrSf9t4BYTTP4qLujIgYQfX3q3D8OQoViimF8VI6DTnR9C1dEsD/dhHjxgUaRaKaYJwn7zM
Xx9SxtLeEmas/wasAscwY0T8iEkz+3aioLs53nkAAETEcpQzIIAJwvK4g1xJ1y+p2a7b1tmE3zOP
qWV4fjC5CZtKDfjEHutuxVhzhlXlQj1GtKFknLywIsWg9OTe4dMzizb9Xg3Qdqk9rLB6MA6AzsTH
sfbACovZpvblfE+j6fwZGjRwUQ60T9slZohW159fOC1x/eDQnCk6HFkCVopRfyMHBKt+V9QIe3WV
fPHZqv8JrbaEGFLu054a3AguUapO0G+X/sLy//q/PokvK91AQp0+oNKiDQCOSyuoevXBp6jQcdg0
niH+ywQIr3PpuKhOQrcxrrp5JVumLAdodmcWSI/J9/KikylnIwgEpsnPV6lKpuMecnwY7wCsK8s6
A+yWiiDcWFDM1ewczPvUck7LbjK7Uybs0GTqp6Kylcxs8ZSTlCLD8hFsXySNfch4zTEQ4mJ6L0vR
i6622ql6DFDSqzKiGpPw03zNZp+0VamJ4kCi2j9Vw86RXzb+fyU388G40X0SfilpHwMy9eC2QPjE
hQZcdRSOZmbA+a9daREhB6KhRdrfiGb36XdjnGyJ7D7n4GRwWU1CZbThO+RWZ3x3O1j5XvdNU0g3
5cpwHbS6YZeCbZtI19qn965YeYEMa5HUkwmzMPeCWCCxOe+/3b/TSaffsqNiGgYpXZhTj39bpcrf
Bg60PgADWLk6Kx3RYta46qLZIyuUjBzEyNr/1Ogh3Bm4GMtb0rd/YwKk6N8HNvQntN36NoE9OEtF
AYmoL/VOMKhvLxgjMQEa58xCc0GxCEiCJ64lc3+hOOV7H8pYR9s++osjioOYmyvR9WgHGyhTD+Do
Uymb8gHfHRH+u8gLPSVhXg4aqOpTigGxzPzAahGc6YovFfh1TCDsNdY6Nvb+HNd6Zc8qts0mJ9q7
u9mxtMqsltEFZF2dxz76NB9cexBvgWgsvk6kbWtIOn43piFHhAvj7AnTPy/mk1TmEmjYTds18AbL
xHu5YBDUpfbq9h+5xNVBZvIhYXvSzf0gpQYSeo30HREZIuAzUCK30hs/uBdKgaZtDLFF5psi5rW8
Uqco6HMa0atKKIkAUVSg9u15C31KbHm1FMy665zLKQ1ZO8nso9LR7Sj0GhJ6OuwXNcOyVdPBcZ98
q7qEM/bBkXk2Uf0LNiewwlOvG5GDx+TvsnLpuhO7ismZa1QyN8mvFyHtf18oa1pzNSXpFfHvZqUv
6zk4lMePD4FMeGsbQgLmdFkF7S3vE/TGp+fjLWUJnrk8WPOL9cRNNz5/iP2vqQi3HLifDEfoKteq
ZI15/8E+6Kc7uf2XBVCzwS9gzU03ii31hoGXovbuQGcQg1M/WK0Mq7H8ilBPMvYp00c5sXhFlqa9
xbYB/+3MGqmY/uDpPSvB6f/ENSqTlMC80ReRF/h/FlJ5R+4s87Y7v7QYgiFD8HlNYtVr42ZocRcJ
6H/sz/VZgFlPJiPsJTQmO2Wdpa0O7M6Xf4+SZR7jPjEiCjFqNBJOl6mzXzYm7L5tA1mr7dxhgWsX
Qn+PXNkBXfx83++u/SAH6X1j42CSwIVwRltybdJKOdGd81R4mL0h6+OE5OeUbhFmHjq8RMCNPJO7
tzgH3mqTtIcyjYJ06xtEMNps+uUuV/k8z1WMjh2r9lC+ZylSRlfKELGHIEY13ALv/Pw5AhS3EMiM
42nyu0BhIJWSkzFe/AFkfAzRBsclCKy1LGk6YyT65j8GHQiLY4G0hX4IHWYKOrBQNGqzwQDwJEBi
xoez58VNEnAjENn8L+k2FCu1ty2kgDIg9tlo36sbqrcwNMDX3Ynq6hOSAlWMzwI3z3gb22F2uxCW
bnKp+a1Y4Ak4WgFehtPpOptMdQyhNh+2dZHnJbjyKo6aHBobiIIXA+4Jxv4tt5h5IRB0UGtZOLjb
ED2lB0su3aTbANtCXs9GrtHT+hrHW/DCF95vlG98LK5t4pZmsHcIgvF5hpKR/5/gmKqaBHAJgC4r
5fbXIr+19jJ5C25Qzp9QaZ3YcdyWf0yixx87tTTviCehCiL0v/Rv3KtKde4nwX+4PPxVjVXy/5xc
NXq7IR8vEBbqmFqpEQWskd5PEJ2KGcR77XkVN5PEXdznB/32zi8j0xXJz/0CUuY1Bahm4Iew9f/m
UnugMkPl+fzHk7V2AdTD/0jYV2ZZ7qL3MygsGhiJs87CTcLsIhhwLHzQTiaE/GNbjuLfWnAhmcn3
+BkwdM/xNQd+Q13lNK6j0pt8As43S07tYO561CltBYiDFyvR26e12StEtVWnlqL5jsIF3P7YEtgV
37MDc0IHzKRwyVY9lDMnUTcxlzIuDbaZvoZ1U+K74NQKTObMIjQ3fCR2WuuxTeTBCahWiQblYWM3
cyiITmPnreO2FZUmmyYSgXjsIe/uuRUyyTZUuONDcGrmA2IDiTBIXXCZ6nLipxaICdLHhI9Vqdbq
oHjh7y6/z+1ym1ytgXu4Bcm0M4qcQID8ppTUwmfHMtGgUFdkAqUm2GGy99DJdo5OFSm5fkHpOM/N
56VIygNL7G5xDzlvv22AJznRlYtRokp2TZYLQeQnKt0j2VL+VOXeyK+oZrJXLpMDmzaKWVZ57pm3
2zOFhrkwFH057UJp8smGFoBLPyQRSzqT2kD0k4wRU/rKoYRFSnd8Iow05bu9LcqNkLtND0ZN3cbv
fJUWTCUdkTqYNKENyL2A5SZbdydm2lIlnFDscdvcWkSgpukuXgMebszcPMQnXRaRIvc94lpH0SmV
GOPTKGl7I+YUHjL01NepfDN17LjQiwBYLeOhONNdZTPEiQnEE1DEfiS9jxzvJxiZ7KorxnzYFlFR
RwG2qGnrPRSxpdji/xnRvhs9Nyw7FBObEGtuoa9IXZ8kNC3441nb7n6MTgCWpd9PFM18iNMfraw0
sAxK9ifTshpy67odlkUnXouGXoQ97/svBv/h4+D1CNjts7SVudhDHDOm42NKIPFi6o23yKgp4ZqW
pIT1LnAL24L3DMtLTIPTdPL+acwz3WBmOu7Yxx14E/21WkUjafuMA0r57Z4QgP3kMIrCm9nlp9U2
ElARRJ3I/fBKtroYl13mY/Plbe7cBhsbVbl6Qpu2Z9bTakbNDdBASCVxpWA/iIq2FIB7/GTIlz6w
IenRuYh62eMavL5XTrr60HmLlmL/Ne5q48iZtPpgnqHPqod1PIxjuK3rs/PSJuFvfH/VPsbDO2Hu
vfiuuX1jap0pdTFW4y9nDH26qa+xZO3xud56DV6LERMSNAd9LbHPzcISzB03nNBSGfPV3PS6rDZG
1IPz6kn3uuDoCVfnr0vULlEqI6e7Chhyv6rSKKUVa4cm3vZCO6Kqsnl48oCHFUkJJRMwiO0tBOfS
UrJoQFVgzgOC1Vxy5/jYNhslaxhdolmUTg5XyxxltgFBirfv+PccVptyZCGz5f/z/zHxKssjRlZU
N0JXTYkVpJb7DdApCLIxFyvC8FXgKOQjuO4B3cktrjj40d7hRozdy3kfD3B5BwXk/s9Fwl2dgEks
82F2EmjgRoZb8w7vW5/wt+bDFLx0svIB9vyf2639NHLz/BsxaHpKoJhwXH+n1JGP7YoBI8xl9Nle
ZR2vJBJhs6MQ787E2y7zB/yxHU7MxWWekf2Wn/yHpLal8q8jmdYe21uTJvc6vqRxUTXFPzRl2VAx
HscCjR8/KXysJHLkMpPwqBydcEOV3u+OXwJGKIRkTFNREUa6M14cDDVOv+ufzVr2HOsVQo99L3FF
yl1ZWsgMWPuRxCOA5kaD0speVVh5IYXtaVFwcY1fJasC97dFSSeTYNWFVrUbkNhnVpB93Xdra7pN
4gPZXpPgUr15yTN9k6d/QmUrAMaehXz5rE9LY7XoiLTm8NzN0LKhpVR/uV5exMiT5wH70qlX51XS
mSgvBh3DAqVmUMjwhthJgDWJeUlxRJFcP9/t3MZoPReZo7n2eeOipib0Xid+hLXHnyWTKbEvs1g9
SD8XTrIPooxFXBPyC8xmVM6mZa0C6/GxDn8iEdwiOr8w2bg7/jmdT2ou24VKEWmhjo3pEnEIwWqR
QHQnb5GWg+jv1yeynyXYtFNDzA5YM284in6uQjX/7SReJhq+u66PtQgdc9joecxcwsrEtPBYIXDx
TImcmfzP0uGQ0ngGgpNzNN3exUgSDlbhLosnA6y6KIIUhFc6egeWK0ewc0bmPbNR5x2FXYEueqQd
YI+M26cHDNaYeNV1D2A0amUKo/Mhr6H1CaIGST4kUDo5o+ObfIDb0NyD/h0oxXuzL8sDNxSeS210
CsKfgQ2fR5MYi+e3y7CbPocxDQhSnGefRqS6lr1mfZcuy10wT1DsQLgtyr6t1iIRx3gXEnEWivuN
V+FaImnRj3ljkhgwVlY6UdvRUSl5WtK+vGJDatgRZn0TPzogErKa3iVs7fA5JFpXPJNDJ3HwHUhW
4DVwDREbuVDWwySV89SgimckIpzGzdxye24EdRG6CU0ihcEvv8kDxi8f1XQZH8ii8JPtorIqKE6b
O/RsJghCs3OtVnnQl7F/9ZddiFQyLIT++oR3+RSkZFUhNGQ9LiuRJNm3gwF4xMJvPsNdcU3LmXe+
5+iUmoNhelHdpRW1sTypDQ4V180uI+RbCXhENJ72kwZrgJvU/NUjwAiE9Ro3/zAIOuk+wz1v5hLB
CPNNIf79/MDjSpctPulAO3gzXJ6wIi3s8/+mXbq5e4eBgqYA3jC7+jNbSAhBnQa04TVDwmRoqTC0
cpzoNF2hmnF+SOM5oSp9zvTBL9026L5r5/In5pm7d8xV9oTk10lxN9XjmxeOWILSSR3llemoVpp9
aM7iwhM2pCOzZgzTfKLAxJ5j0Q5deCoGfFQN9BXEQhT77ErMRKZBl16AGgsmKfqLPcY4BXK0U8gC
w+ZR5yd3Wl5nNbqTsgK5rUVYpKDBHzgbl/Gk05X07F3j+Kv3QRcnQKxtTMYiEzTa2DlTAR/U5sTN
EpCRlje03VJjS79BarBqGBQC7n0q45m+7h1tFmmAAkEDwLYPArZfCVlw5ICCX+WZASz5Dief+/N3
/uKN7rSau1DFtDkzth4PhFTnBn1tbxRz+qBkDzjeIqwRg4T4F4JtE+3lJoZ+/lblpd3DaExzVX6L
lZyfqRM3mZyoMMVcB3Q1k3vwFxrf/8j3UNYxdLzGQCAPcrP9VybZ+VIhepYhM/lg3ezBbdAuqAp2
jd7fpLZxM7kH3+PVPwPyyY+QtVaAYAeVV36nLlhwKFr305BdQ31e5Uyk/x/S1x7q+gyMoNN1y/j9
AjLT0OU5FziYuiwSvFNdZLJD4S9Dc05XRVqNp/GM+zgK4rC2pacM5MLWiHLSJwBpwA082hvCgkZw
fCxpe81qn50KhHVcfIAVY6HnCPOk1X+JVmP+OsCBP6IV97wQaAOiamF9xmufBgHBd+pLVA95N5mF
DF4aaQzBwhMEJkz7mL1YwwqEKaesS4Q485ka1RQ2151wRjKE3bWaH+/0SNZmVRMtTUo1o7E+aVjT
CdqH6zat/tAQ1TwCSEI31Mgey04QPYU5FxiV82vcYeY6R3u53ZPlqdvze+3rbZZIwwHYLAEsxTGX
RnW54BycJNsLndmy5GqsHXVunMtBW37EbkMeXPrAFRAgu/wIDgmz/R7LgCAstx8iT0gxfdJfmEbx
pjUR3EE998izxP3roWUrUCs4zpZXulNINgwMr2Bmcjg6BKW8vRp+wjunEV/7u/AJRlFFazmH4aiH
PUX2fLMsuqTG4RJDCDq7gVnd497XIvQ2AoA9x2q8pyl4Xr7ELy3J2CPnil/S/9d2OB33091uBYPP
/qUNq278GMRqY2Nv7Vrg+RjP8nPdL3uSjixqzZibZIpDSEoZM1Cse6PWUhW/7BLcq9FnLTteCSIs
sR6EtgkWChXr/vNlGDtTmtRdSMtcz1XFg9AxMHxVEzlgVUozqsOmV3mWs+FA4UYa5aJg/uQuBQUt
SvIYxbwbpc+ebnTw4BnMm2bd9eK3GNvSbF0y1wfKATYIXlq7lrCwiYVqeoHvwS48r5TzA/54h0BW
X1iGIswdfIBi9ucRpH5U7Or4J9d5b26DyvyzQZe5CmwbHf93bEJ7lp2A/as6QQfn0CtChrWPZXaB
2z3dWLjfI9AgRS5/kEYiMjVBNIrbsRAC6hwbYTaqyFwkJkjEHWn3LPUHlc0T6i8Za/f5achFtwxX
L990qzt7lVXPmXPWzROtAfTCOQhDx8C87OOC5I9+KbyGKIK2h0rLxTimRBle40qmecNsg0dU28yw
nhT75FTeQOFpo78Kleo5bpJxuew7N9wxgEnccAoWe6/t76DAsGMUtJPvRKxEPinrctO6PjeFbdeM
oKL4MZnFdUAZRUrtMHruj+k6/tzso46Xk9frCTaWalgQfDAuUUw2eJmHwsTD9+fUXiY3pPqHGLS7
2bMBnhY7gVcTsOI5P8/YUNgw/GrUutUK0WpxxG+a5PQhe2eIqE3XbaS7ISy1L5dMqMmPr8mPsUYa
bnM6jxh4Td8kErV47WrgZSbWxzA1uZMVZIK3AVAUcJZitGp4Yl2boGge4CDEv4PcaZX0bUPeWkbm
xCYg/4vluenZ6NZSGGbb6naO53SIt8LKHqTPAo0JZrOpZV1lZLKR/5vlNbx3V4D+vesClhBtaOev
3CUzNnZ72H09nR9xjv8Jl0jCay+V49senaoEYEXk6nCwwWzA3dnmWAMmWaJiarN0h+iSwB9X/4WL
owcjWljElBV6wHJh860eDpwREMYNN5gemuocABce18tpKY3Av+F2y2dG8YgjAKVlGRZAlf5dfPsZ
/A0FmNZuwnRlUpK+uDe8UveeYRON58J4t54PJBmZBJverMiwS/kk8un6d7r/gcH4JfSoJCTjgnl3
DvU0+jvbq9kxKlAVTPkqTy1CWZ7Bg0eIPP2NwffaPcaiSMHc+chjcE/HAYPkEsG+tcp1SkzC/URO
ohSn805WmTlvmD7iPOpG5wO8GdcLHDQu7H7Jyw4A1AXaetpTWL+RW0JJTPoZcv6UKhWGlW0x7PxB
P3Fw4JkqWwJlydTFsRcg+6Au78VrDU5P+4bKy2PIc6UGfXepWTbrnLVGi7wT9iGoP8R57TGR5SVs
U94DPgoVm8+B+CJH/jhWr9P7lHSyCV2Xa35HP911/ShHnbaE1ICPhV60gNdDH6YafgWEAVULNMwH
OKaKogTdgwCdFRYo/f6HXJdLQXU+mgMdi+KqCkb/VgSTaAd5NxWslC0TwUunfd6/KkEcxDBnUUop
qD1lDJsJkT3TUi10DUN0F2nZIIG8lJyl7qazy4tpQOwkJcn4d6ayfFEKwEvlR9m7/LOva+lVms3A
YYqXK0NPTYC+1KScHF34b2irUeXQz3qkiAuzAuJc7jYDOnY5IDqBs1kDLGr1/jQzuj0nE9rHndmP
Fy8psak2FkPZDcluXDa881wXktyffEde0Zi/jgRPjE5SjTFJH5enZ+4TA6EKEGe2UukbzkJZ3UBV
AdhWDhyDAJkCv+4WHEPqp4EmUvGBvuF9lOBEMbYT8WAVxsiu7jKzqywGkIHWNWiXTwbunH+HigO/
BO0mfWatdCQom/zeLvvFaEYm6HiJelVXP27j0RxFEri3MWdy/XAgnrQTrxebWrX6ue1r6eB3PAI2
AiH6qjKo9F7ZtHBxaBte4ECJqBx6TK6r9mgrc33f6U1mF9aR3RItLIacgjM+A1sPWjIgXYZPzaQw
2lY9s9c6Ro6ErAuj9pfuYXzwoP4lOJkVJYbJv6z91+ANyq/DFeaIn6nL+atVbjaaLTnahyGhyAWC
CpIVTrWZEcCdT5aLkR8DAQ4XxI4aOjVqAD+OKEvX+nwTWGW9yCluSrW9uojhOXrzP3d/uQ/UeYN8
pxf6UOdYAc5y/RCj2Vrzk+DJM3fnDmnK8TfYJgRAcCCKcTrBZkySZMDWwkNdHmzswJ1YYc12MCd0
waPTTNqhOttj5EN2v4LX8dX9HlnVJvCD/koP90SOuUlwI7RWq7XiKv1OX+gSRzKN7XXNdUKXDcii
JH/f82b0dJYE/gOvP0BbKKCy5oTBbhFEx+uHX+lUgkQT7Twl49KgVgTyibCQP6zNQa08AGL6E1ZP
DP6h0HKE+W1+OGkteg36bzfh0dnDQ9XkpnbVor6r1stXAc/boMmeOIoX9xw1djQLWDWQ0JXJ2WtH
dkQDVGOYLsvC++qh4MgK6ieKRt/ER3KMDiWobLfJ/3Yl+1PvgNSmNN26EyEpiuwKIxpste2EAuCu
riw1kC+Gqmnmb5yCf5y1ghZjodyqsuZLpSKjHsqGvk6/02xTPFn3QL0C6hTSngFJKVxIgcydVFzS
h9kPasrCsvxBG/PSKVHkThPlO2wCL81NtvFI7H2BFRbQV2PJn4nJzf4AqAJcxOU3vP3UUaud6EM1
0StPI3Srp8Q/kYETT/xJUfOUaLgyFKx7QZ3STXi02GJ0g6aLo3d0bHag8vdaDJP4pfY8nH5gcn1D
uiEeEqlLU39BxpLxLb57oTZ/5yzz0rIPTWqyUuFpWVzu9JrayQbNyzGWU1lDk5GAb8IJTfvTPamm
lg+vjV99miMOihYkgRMdTO5SQtXfWyyOg7PZZBcus27ZCnjZuIraa2FcvuzvO3cAZXyOU9Vufhqd
koA2Tm/BDH7BTH5Nl68tpS+7CgKC+8LypkJeglqNKO3BbeCPz/mhSWBSOOFHVOYysmT3MlopYItx
w6lo2mG+mun9TVIXgWABYm7OXY7g6MUdeY58hLaTySBW5iq+rFs7/S/ps2v++KJi1HTI90F+JWGO
N4zmg9gJKnlTn6AUBV0OasNVQLjib58J05u2ORSGOJOcRMOQiczNlwf45Ipl+QcFnx8bbE0TBkBc
nooVu5rmKMPbhNHyAhrNCbrHLHrdVwrleFkkYszhGRJgDPcboalIlNW1lNSzrpIgKyWeUztMSZBm
Hn7VpJKxsFDeJTMylXoL2UMyJafH6znZNBOYv7uqiEPFkvy7h+LfhvMVXnD1N4IZRNg/Tm/oUeo/
C/lTbpiZ2mkmFZ/YwBIErzYPHWuJDmvKR7e8ysTbvc/GqPMU19+D7DbLaCfDQPJVb4Y2qFYWmMJ7
bRonZeRGz1Z9KjrgUxDf+rVmfIlogn71Iq2PK3pVSBFLrkHtr+WMF5fRy7GWG0bw54+RL9Scwrx7
jfe70cL5PzrUtbsWZ/pnbV1bAFP5AC+QsNkBBT2cMfTPMk11SIfH7lReEZoUAndqhZocbjUNlxRH
JQMe4eaUE4gdZGOuKTE7ajeDKbwqzOKTpMBZdl7iO6I9uxdjkV6VxidRYzmh7tTLmxs+QkxSnfKT
bxDWhZ/UAs4Dq7++4WDSusZX7t78w5hhBjD/X790/cQYBCm+/E88T3KOtVmQSRSsqm+VTXB4URec
l8bX/PV6ui315yr9hnNhCNF3Ed/YrprxGI/I90ZTeipD0Wm5zGe3YwBaN8kp+2rRKO8cidVlswNg
gTl/YqNq0MMmkb89sjeJDljPR/5WQrOl7h6LtLWbr1yRpU9S9exsut4F/dFtaKWM1gUNxy08J6r0
oh1BdnUWBJz46r866Kyo5Xoy3X6k2Gs1Sgj3fSyuXRz/vxgRtyx/WxBwdOfl98iaZ73bmjL4wEQx
JDjtoBV5z3HUKeM+V1b606EpORB/qMJf+/xAhW214noA2PnGPexMKQqRagHrEUV2QzPN5Fhbe0LZ
m9O6W7fBnLyOoTv6+fI5+RZ3nmxjhbveX5TuQmFtcqk8g+R4Jt3TlJz0CTDpS4YtM5umM5QVVvEQ
QILMt8XR4ZDv7C6bWNd84D6Ep56759NubIHq7NdhFjPxfuBUT3RLXVJKURcnHwNWZQv66wWPfbHL
/shFCQVfq3pfmW65HqIuKSD/uuGNjbS8QVLB5GuWcimFS8t/wbXCU3zqAKpQ2CWz+YcJSEKGecUW
ME4QPF9o1ekrCBbxRFA/8mC9H5NT43/rGO6LRsDuLX9v5qXmVbrmXW1NmIxFGDxIWxV5xrKngCNh
iHwRJ3XMopBYcYmfpiXQck5RTWPJka/KFwEGoR6UsK2+IWvl4JDEi+nvF5kn1dmnGz/lmFPcr8uE
2jUka4cvQ/TQXjlCay1bsA/iDkrQvD2UfbbAbintS7baPyBYFdQV1Lwo25/RmDfeez8+W7rIoQOd
Xo57/SVskAOVPOekIbhOwfKLNcNhTKtBjPCCxK18MSciQ5CQoImdQNvuzs/MplvB4Xk5CPz+7mLq
LJYVu6BnRdCTz5mVNar5M166mL3qaOaFkPU8YtYVGdiTbhPJGE/yt4ilArWcRSTMVfcpVuwcBYg9
MGt9mjUXEBbeNquj3WcIfeFLgkMv50ItP2yHb7ON/p6zqVqeSoYKUw6FbW0NiUGVZDezz1BJsi7w
bs23Y4P0q9EEWo3LE2Kq7og5qW72wR+VFe1Sgck08zSCNbzuuOqvUrFLN3lps8YA7AqN/qXdqeCH
jfMxVrFmPU1Ryxa+Kf2x/gThoXdpn1Vz6oefZxxV1LNFZ+cQnRjhSWLuP0lEmkKkSgaLiAeFvN22
jikqtWf3qqWo0UDFWVs4H8QeSTo3xPBol/mLMB3CXsLj0E57mlGAHQ1ne9pkgePCTFEsgLYx8Wq1
SGJDl55ctPxcrAkPeHBga2y1otWncJ+xJHm2U1rHU8pVoid0LW2qyk48Q+qyKXAiOvMiBi0Ek9Bu
Vxs72+7PcQXB+SqDEqvjatojiftUHnOlsLaxwY0u0Svc4nVcdwTnZd4LAcxkUvnSB8bzvOMXS9w6
gRtQHORWkXbQsVopzayyic2wffF4K+IE5R1j1LU4bxhdyyfgga3LSQSgpAO2XHaWqjGqRXCQev4i
IaNFpT2rq3lyZtsNGD2/lWH9hIQpQbHPWhc5lJ6EF9vGU5q/Qbl43ekBkvoOtJp6+IH2IPMD/XNS
Rv8p1kSV1igtHICr36S3HZlKNr/N2Sf4XgPUeU7y5x67dk/EIJjJYiLFiY3bSS6fJvPPUNv2Le1O
DFggS2UiSd4+zAlD3q13XnfAZbzTszYw8cxnTgk0Hn2EeG9x91gP+Ruc0JmllkRz2nEDSb9FMt/t
qJwDdkfiB8Zh0NhH2LVO8Z9/MKGrpnuCs0dWLfQtKL2XYjPEgZjZliO69pQxUpimY8AUT82J/gK1
v/UikQTGkAeGHloM3zVQ+tgYJXrT3hGKg7STQ4l/4qJQ/IEIwTgEAuLtbsalAqAvs5rqveSJang4
80tZklIhqyE/VGTjlXjlG7etka0hFLqFDPi5vbB6UVkgnv2CwkJhoJeJJtKGcuxVZx2/JsMg3wx/
pDWxII/Z8UoHvhOYCLX0QukMxJuxQthb0LOF6MHUzFTUw9uP/lWtB4/V7boM9QJCS5aVAhs22iy7
6nFqkZMkgjdIzs4cbdd136sCNgAEe7YqtaDjXZDXyJb4UB/EY+7dis2SW8XhhkZEZHuZHnyuwfp1
kTgueiuLEv/dpLaQJ5BFKe1vSgBkCVK+WXaikzggVaTYHQQj6MtTkfzMg0G9u2TYxyD1kIRwjzqz
1tTFq6ShdK6PFXvOQD5BlfB0OUU8Yh/uqebS3ofdYlj91JZIo5IgkfBpikjsq94fbtEPAIA/jJie
ZJpL6y+NKIq768eOBiZfNkZ/sTVR3C+y38620VTh2gzD7OR7qBmOwWoVPjgfiVqACAp+E2IryF17
QZ2L7ZgXvoFRXvHKCJAd4guR9bEJ+nvboDlryiTmt9/RGdSMAWeHb5IvJD5M+NgcOUrI74pPcsBv
N0L2wawoRMwxJG4EvL3V8ktTEoHYUWUEJNBG3SJZnYwtjaCZYBJMWagkWNyM5PBM87vaShsWYRjK
qS/RES0zPDx7TFfok0uURF2XC4AHd7MXDje2nGfFr6revJ1UliydPqPgOj8vLD7zVqLpu2m4CoeZ
jMS95ZOekqHOxFKS3Q8C9e/um+dod1YDSsIF0qTFljDYRbwG0JTulq79yl+TJz7/5fnCaIyevKVB
Qw2xsoikPB6ZdKRkGV2gMS13uQYuq2L1qSfjGzUInfDipzW7mqZtR9IIQn12bdHmi/j6LRLINwsZ
oWXSsBkmbRykOaXevMOjWfRLIF6zKLery1B9icBp+KnuVZ3TUY2rJcqANYIMHcys8z28dkQUXWlS
YyJN2Xhb+HAoMt1kFI7SlWDGmWZ2vB6lJxe9zx2KBe7F168g8+AQr7nBckLsNWUkjGyDRYbXNsge
XpKJ18TtRbuEoJtuYKkYwmxuJGHbY8RsfhyDaV0vZRm9lOmCN0CPCpQcHAKFFpNFl27qOthBGtbr
M6m5endqmLr2XOvDirL/6PC+rnFbwwwt7NWiJM5eH7gdJgzW506Qb1K0/d+Gfp+OsHIRpHQb3lxo
LcQc7UlMqXzBX97DG7Ijh0bchpqYgN4q+jBHePlEVLHBYuZfyQ/2PkcoAwhc3WUCXgomOglFW1oV
BCbZGGGyJyq/2ZdsMN0ZjSYtCZMW6qyfKEZqXbc9oyTtWrhhjwYETfelV8oenX2Yrxbn8GOozptm
vzVJNGxpVreDlaYM/wpRxo4EQv4S2q5e1shpJUZqxbl4Bd3bN82nbL1vXWdcgBS02vbklUU8L1zc
Repch5TjDNdoRDE8zH4FlJDfhFD8aouo3gBHK/PTyK4SjH9lXbqzyWRHIxfeJ7NVcFtsrF/SZLF1
X2IT3l4CHvWlFRrxQwNo39qFlIu2AqetQQi/0RtEL3ouNODsUJNouy4OJ/oL8xKhVYDOUcorv9Re
jKB92RZqhwojSa91Ww30W4gxAjSUZuJPbwAsyURRhHxOg5d1v2Y73VXMA/VxBWc0XqG4yEZRHQWu
NIew9J4no8TWlMeFWXhfiK6/q1w5EYNSl0k3Vwy4SaBv9rnZKP15ZsXPbs6QwAWzQ+XFqSajJX2t
Rd95Rgx2lNxAm6J4bI3cKyFqa+DbVIe9h5sespgi1h20UoZ0MWPpEvaAE7xxsp/tO8cmsJH1U/Ro
azZGxZJwkV1omtggmRumZ7Y4CmKBqNe1oRx1VxVwalCCKfb7xaiu+mKKLKlukmE8RS40iy1plEUx
HCV13JBENFSSKDl9UN7hQrR21NAMTKPRcFUOuKqc2ftjqyodOe3C3X8taxqFqZvrODOBqlOmeD8h
OYSRC4LMoyew5M27V4Vdsz7zvA+DYiOcZDkMao4kY8J3RBkDnTq8h8Ex6wSZdsytJGTg5EW1A7xo
PRAUvGBXJbjzPFevmXUgBapSTH7Si28wDmGkDz8mjsXymwfJv79me2DCDKYwAOkksW9bRehdEEKl
omTjnPayZ9PtXKhdzpF2EN0o35oW7aJtZhsAtGtq9U9+PZWvJp/9LtXCkMl7Loa5lKyRkhMG1eOX
nOFyEjJua8LvXYHzQbua8XcdzQbJ8NTwWpWG/G0sPxF4/qndp7Qk/S56z9ZjFw0NzHmtRYRK4NCV
668SEy9pLLvR4DDPw4UqulWxEC9ZQNDez+w7kMAmOUmkrjgnVULqjitds6mvGX1OCbpem9xn+poK
u9u/80s9mL0MDKiti5eX9y3TtjaJu3Ch3c/Jh+oiH5uD0SxWQXw6UG3yxISpPC2SIOBBeh6P9yrO
YstUiFWfsKKmFuIzTHEX2VmgvQ3SiBQnk57osiFeLsjXJQaWfZMRiuaf5FFKqjAo6pUWRNNgZZI7
GBW9N2Drx7Yz52eCclf7Ex1rqiNCQqhEmapW/rVxVeKde5CloXXKwewARQ34nf/9SKVYlrMvDGG+
Xhu5c+szi8iCpycki4GVYiNSFEwfLjignjuX0IrVexJ/16oHCfWM0yiZM5Bk76HaCKzfLlzqflj1
ssccfjOdCmtj+Zn4XzywjgMrC8gPPqtjLiL2pU/Fy1wbZsEJnvi6GoVKcyNWSfCxQ9eKE/42bELT
Rj8bWASK6dnzpFuETh9AT4M/8gOJ0x6IkNvkM7RCNkRB6mMhCFd4egXarFP0vxmnmSeT+m1LJqXX
tyc1agb/hJtQpBDIVL57ASifs3OF0jkQ5IaPAH5fh6wyOaJ7g/SAuHWxIq2DpygW/t8x0sxeDAqb
VVjqXvZLQs7SP3fIibU8Njqteg2fayptDmeJEb0iWImQHl9fQ5x7iHvMJfdhxVlSDz7vtVHZman2
kBe3xyirAUiTvKhAdrxhZTR7YHURRvEInAOPBxHTMiqFgo9fXx7itHXZFZsviLI7EJgiLs0R+dbE
9qV0mZTQVWkAnqrb/2X9CZvURiTiGQeVrVWJRAthY022ED+D8j3zmFVgJCBQW+/CNlITXxqyEODF
gGA2m3J02P/xxtM+LK2HOQtxppzHbGg8zOjSuMg6JhbGV7ym9t/Iw3dolcHm+55+sYd7ZDsW+VTa
m4PqXZQedDo0W+UtiN92qcsBIxqbdGBcOHQ9GEc5xRx2ld0rEAAW2PbFQyCLU1jPOhTnwutcqg5Z
v24x2y5o34Z9yh2ev1qXM6i1UaRt3K3UCE0MSof/hRKGoTCQMPw17q5ZPyZqopZSM3EFnWo2GrQn
S9LqpORgmbuBzco+F9ZL/0v9Ez0F0L+BBB0Q1S/GTP5Sy3g2VW+7xw1AvflyswAyNIaiP3jaRYOc
7WLWvpZry3Gq76lo8dPuKftaRTVyK+3OWHHQPgg2hVQ+RQuKrGfhKSxcuLIecZl1XOyhorGCGRXB
Iw+bxqNN6VGwtRlYp91QjUzggnK8gBzpkYIYFuJdhyE2NNI0xXTNsVBCVtFpoZDKnliYgY1j4/Rz
GO9pz9xKsIa18EaOZ+Tg6q4JWrTf9wx7DwfS66nZyrviUqI1kUattsJm/NYsdiMGWP+qfQlhkNOr
RmAsuzHXZXUlYm79b2bkq2yqFy66ejbViv3v3qk2bUvTs7tjdlXOXBvDUAH+t1ZcBg+cTTOIo0Q4
fgXWtWQ+SMcYLsphvqEYSrj9m4pRsRECtAWSTEQNpuVH9NtRVaQ1vPQncVJtZOF1S+0M7ak+7zer
stCpc3EThfUYyOWL7eyQGrCA7d4RXKCv9+sVJGjpEhrp8IBQGM/4pFi90PqseGr9Ys/zUMxtYY8x
XZWf3zx1eDWc+gJqxd4cz0o2EJ7QJqKUUuNj88GWRZtkfPXR+b+kdueepEn+cLNNOPWOT1VCvD2M
1OAe16XkDHrtIHdL3s2POPK5euCxhCB32e0sD8/dryWAfhMAwEcngFlNlvH1PJugcvJw/jjlOVJk
bvy757yuhys8cheVj1KaIK34TzO1Ee8Mr9O6nAgZb9kKteccUTtELFdpUUC7N1+qUoX8dhOi02aH
kQZJU2TaiDH4H0NvnOyaV46XCRrSIBjpOzptGEN8LT0mA6l4XjNFDjiQIilruAMnf42ZX4ynAEMs
3PZ/KMIh5eEGv9eODqm+KNmlnRVKLNihi661PomWQ3d9lgiZvVyjYgnLOc4W1iV3L/QLWSJlET7d
9Xy4M6UnK3YB9WI0XLc6BKrxwE702rheVOjeSvIGMFJsNzUsCXvUR3akSBneaBIj9JlCIcKW7ec/
j86lbCc00fnUO7R19kXnzpdy/m00FK4BwbngwX8HcI83gTxR2WNt5FD+NwtN/sHXVAecviIdp3Gj
b8ga289a3YWHnS/nu5D2Yb/ngWl0cXrenK5pdg6nnTPGxqIyMGeY/fgbfmqyBfSW3B2bZcrVZS1V
xEb/uLOEFF3a1Z/UJUSXf+Z+YVSajts9gpG/qmDT/kPacukuw2muLlzDOWlKuh+evjj6dYOflJ7X
OL4HaYKvm2DikxahRwtnD5OuyttSi9y3bWR3LK6EwP+NSwM5andyXOrbMUA7nRpgBLTN4cErF7Pi
+p74ZGrjMqcYJvWVR30N8+sxqMk34nZ4P0WhXYTpA5JUYijpx0fV/6nn8DIdPfhdLBenm5+XbjPt
2kh8xJ0fTPUCAv/Rclemta8F9GqjVzYGQnYASVQvNIpEciWu7od2xTG9ZsKKlfobKT4wXQy+qhIR
zX1wOGAh47vJnv7dWqXrbKeIYOIeo3HoOYQtWSqrXh5lafJGXqbVCuZuCMZbX5wcRS1+lyIskV0d
l1K5vAR4KWVbCgWeaash9+a5e/7bNu+099WIIV0qa2AzrHlxjemo/3jtruHDtnnYb3SssbiTna31
Ay+8Sg69nTsJFwe7QlMFu/Alp3Nw3tVXIJvxaLgUby8uDsWxKXzucXgG66S9ycZwG7HzgYroPRKk
JCwOt+DJJKsWobNUsoMAF5GXexLGqkdrfvnmC7VqEQVud/tDpfK5ScqjFvcZ4s0pJQRW3iAZeySR
Q7BYZL8B+WE4bSl5T2PjXrUUJyLFIsz0Mw1eelS4FbdERdMoULfpxeDGbytphPoS9+2iKdBCS398
Rq9xh92DVYMZB+ySMINEwpzq++63o3oa3zoZk05EN3Zjh92s3P+2W4+dAoCxviwTFUDCwD0mZf4R
vDkGg5/5X32x0q2HcaTx8ysloc0I7ySHoRsBY1HaZ9aDF9flQsMoINpBR3xuff0dIgctefQzaGso
uOqJr7vUTVpJuS23QObQfAViZmIqdS8OQO3L4nTg7eVXIwMldFV2o2UpuUi4UBn2xLsCvisDLGeS
sUiIiRgwLa3BYun8Q/qEdlD0isTtDGTmH/VjlrfDWADwPz/iWOffkSHKwsP5Kk3SivAg57P2GfCU
uQADvQYqq7l2iVuH7sDgVLrpsQeyzfL0bW9QVz53yiMdeNbF22O2lHypfoqoAk2TB2DQiCZ7JTc0
INEArt1AV5CcUe5OL9tFf8w3aiB7I56G0xQ2IT2jotTt8JsrJP0ugZqnTVIRmSnR4gclxyTxs6Oh
L6WxHDmYaRn0uF4fPW9V5jR0LHWXNI39Rx3xuxTdJchiKJLBh+o9E3SglSFAs/v9/xxpvUgPt18c
fN7f40QIUXIeEjK/NJUVvmjdm5m0Q1eKRB7rUqHS3rtLncCnt/L1I7v6tAH1pDVdGYIJU+CvL0tt
ibB9g/gTMCdsmyEmBFOXSzW9WzFAjZjokPZR3HBExS02OHXt/QsZlRVKOThGtK5Y1BTAiK7QkU2q
vccZvM90li9zp9JqiUgTGeBo+tBtmM0FB3DfKU0ZWg4lINPjgwmht5/565h2eCi/vWxMJRPKmu2S
N6pVHz6wV0Vahn4ctAIE88aWufw59N6HH8UzoOeWXfRjyTAm5ADP5vqSlIihRez4S6o9QZR+NszM
sVaujH2pQ/aqru3mX5qa3JY9Xfzt8l3WpYcLPeUysYuRZwY6pKvGJzGsfRScVbtrAyekH95bLSEU
2JeBdqoYwdHFmxFusbwsyBwvJ/IvYdC/oP14o4NwIDISeSPoRHeMmmafbtyyNdJwDsmLikYlZEo9
5XVimBQgOkuziCGxAAfR40p20bITeRaRh5xBHndnGKD/EmdMmhcYNgDLQcFmt9luC2uJbSTYJzC6
omRx/1TCaBcfRf8cGs3EGOQCYDYQb1nVpompymkuMILWOphLhyEVP1IUZPhagY+umKaUCY2044WB
AFEOjyBoSnrFe59UlUB7EFXxQGSHkcg0LKzbmUdBakeuRX9D6AxhrsnFVcxyc1/LX8XkZDr/7xRE
xZgKf7Pp354887Fc+vsxuKFL1OeoS53iRviT4T9vnXrZZmjF6yZLucYnAjzdW42HSAYF7LyeUK1b
iBoqSlKF+mrFEeDS4qRbylg8MOHGyDm9q4QN1uRhJ6pL9l+wc58vet3ki06U4WWI98t04j0BdMY2
4mnpvx3QXnCq2niou/bZgowg2fwj7ObHeY4elSIt2QtV8/Xxq+3uXf8qX+iFJ6y/BplNoVwTxqQb
0h8ETXQXEqRrPBW2FtmAdF2LT4TDdg3waPIV4cpTljjLj5Y3B6nHePx0EsFAk0+6UCI1CEyDbTZt
wwrh7iypkjc3/+3hpqPciiu9PWZs2xmOeOjcUDLpu1ARhR6ov4CZyrd1S0pyJiC6cnev0SMUhC3L
mhpu8clcw6aXdzq6iQEXdYCTsVt59++J8DohSOsq8Bl/DhYqEdczL19+CQYnN9688qrDvDl7we82
dXJ81kc1zyn+lOgkGAB3kUys66dbTiwfujsIUs9u35bRh0LS8CfW6saz90lrAVQN0zA2BOACL3Jn
c4VdUWgppzkQfFBZrJNMNWN02595rqzum8DcnlbOAeZSDqmja9TUaC31wYudcT31+KXT+fLJWKCe
IFXY4YIRNwUtYlWFt5mzso1GPz+mdrx18QbCyI7UUf0vmOTqDYNxDtAFvWZ0Raw+1oElwRMD4XCw
SzIbn/R130ALZO5OcxRFINF6OjxYo21uwDvSDFLfquvN+XFlm/GLbBYbCURmBbreHF/qTkBsV1Sg
40Yw07s3I52RreUd7Yw3FRMNLWHVMrCvir6nEi5zWd2hp/d8rF2aDmNt1waHNmcuI38IXC+tlHl4
D6qcaKjbJff/qZDgEK/kEPW8qhRIqJwU9xS6vdNgZ2hlAYWmC48RMVrJx062BL3JxDUfODNbe37d
PO3g4QAxbLw/uz1DOJTyLBJnFFnCb1pSoe0jAzvImL6ATDruQid4+BQ3gMhh/sGz79JTXfIVMmQ1
SWogHT9DpnPzmh9uMTl4QgtH8JtqQ6+IysqV+JuRd6dELlKUlGF0c/QV2BVb2dDn+mLMhZfCKMVA
qF3zpNnzTxGrC7LWCJuWhHtUZKG+2LTXi0YZ2vC15Nf0YoQM5tpULqTG7T4ziFa2RM0cMjb83m03
10LCNYaTG0M28pVpInBEGEvdWCwkbS08Qeoy72UiGhVQuYQxeuQWqBwoAkGhOpayE9AUhfZdAb6X
qnHwEcMTdbS8trK4MNZvHv12pJNJIqoQdhNXogRvv/EMhxYCAPqniSr7r3Wkn/O3zLSFJKwq6Fsx
wKuFjMoU6/iaUx/qwGcY4ReIynS3UPI423oh1LE5hjs53mFprQQz5U7FZiKuNGewskWA/SlGCOte
BbFiZFj6qkKZUQDT/0iBJeHkwyVrVF+A6eozksrGopVS/cKJlUNaAtJRTbMeETjnD7sDugz9SwTX
BZVa4VRAdlsU9HHJIp9/3E+pFnC2ninyozIYvnEeVD8O0p0iK48sAJsDOSE2G0Nuvk1f6c497czW
vdGjwoeUnnih/aPk2RZMwkc36uooX34aAjS7iiVAMAX0iYkDIptNQAhcwbnfMqs2cJjuIB7WwRh9
kAjJMkTxUMhNguxzIWWR9+ejaporyd58ZfuNrwer2MemqKMkK0++Rl+SQ3/CaEDV1/0I+tvuKfVW
M3M4Yh9JS02jRJwp0Y6uGNYvx6REV1QXrQCIfyrdu7b21k/cUZsiVihR990lafVPnVbRnlU2Dbwh
AJL/TuI+0rQy8lqwaali+fDK99/8IyZHru6I7ELOejoypiq8Kd6M4E5VO68uqKZORa/oTRpki/aZ
Gc/NpZi6gVx2wNkoUVYrJAVBRYtPLZXEmnDEZXi5zSaX/Ee981+pKYbDMyBya35HKeITR+vPBPw0
WQKyzEiRo0A8D0o02G3FAh6hRwwYVPbtnUrz8vch5G5i7d77XNJV8eAR8n5ikNpTH9Rkqa3RJKJ2
KY1OXeNCNJ1MmR36t3EgUPFFHoC6RNA4Z5ivNUuXqOZu+iVXawE5FetNPbmGIVhJ7lQi5aiUE2H0
XfTsmU76V4ox2zdDmNs1yAKYl8SkiLrcqHtvMOIFzvCeeKm1U8Br0Wgg4UrznyBQwUsIvELh2/J7
006nv/7J/4J9ykQ3V85jkctjv2Sa0aMnUl4Z3GtzaJp25auebK9KIErBHzcbaj/ewF9/f2BhvTTB
am7oka9dRf1EZyuI0J8Nox3lSs1458dJOEBbAnCVgmIwkDKRRuAuHhKLlY2d5VuTkcCL76fxBeK8
08xwbcVkb8CvBdL9X4+dVWv0hPWhS2aeug+g8FGLzOjFFefkzH/3XxI77QEsDfMpBIl0wuZbyKi9
hF9RwQyL05/hJLAjkhnuHhxvp9za8vxoz0JI3GyR2C25OGhHjJiAgNUSaMVf6j4yC1jYTZ35HOJA
JTq87EPYQ/8aMTXAuzjmdGqvzhHLLLs2K4QfI6DitHmme4axzE4moLxJBIEKO+YSPCLQIDliEtBR
eUcxuSoLBH4WImRsVzE+Bvzc1NIt6ihCPndjGZzFId4DMZf5buaIEXLbRFyMTEFk5efxMnKFHmfF
GfYGAjtu4NkOLk1tsm8AQyHfdGDASKNd1iJbbR7DRcD4G599Z2YBP+Jd6UFk2wI/osIubC9BDqH7
c/833+MDxUaYaouj16ODitb0pNHxmK0MmKOwr9Qs8vt+fFZ6xZypPZ+2ouEc2baGC+yOZ9ki+fXh
8byhLs7B4wIJFOkw7dXKA9eXGNPLYAQUstk6J67XONnjANO6mivzQlgOq39V9+L57Xdh1WYofDBk
oLo79ztnAMdN04rw1l+hQZ5IuzwBjA0n6YsIUWbcEAhuEAc5xjirFs5m5WgF5MvKMUg++xXmFPBR
NZ231tX86uoJNMMhOcCeLEiof1fsQCH+wolgGZnvwDRdBLDCbiXSvuHExdH2QSm8nXaRuDE73Xui
NYQZ2CUz69CAM36C/pBhViceKlfP/ksiPjzFScRt+JpwXkhQ1H9xPuq5F1bVtuj+sw0ggZjxtIYN
M0jzsz8T6VbwpzmLQUYpSt2aixbUgVMJkukT6V6qY0p+Yw7ixe04+PyDpRgAhVdWcV2un46PECwT
ChSYiia7vhYHExq5FmaLWOfP8TI9G4/gGSzBy5BUZvOeP+2AAUc25h3XbgPYDoOEqqmCrU0tuZyU
b3WAWZyVE9wXeRFVRZbc+dM8KoIQ4tjD0CxbIkcVtObqa3Vgw36YKkqgYL8+InxLpjBrCcybC1K0
49Iw9tnNfweJvd+Js16oVrIOZFZfmi7FcCepFy5MhSGFrG9/93JLj1aS1cT00ttU/6+iBvVi682c
U+67rDm/bjg+WViVW68kLvs0uuvLwbW70gX/mmY61Aycsr4BDvy2oQhcLXkI0Gv534LuVDSORvxC
SvLW+/6NtrvjmV9vYz+Atfe+zBJOcqhyjsua4OLtuXjGDX7ARTigeYCoEOakjWEj7nIUfYb17g7E
ao3wkCiAG1jPsFhR11em/uuozO1qP60DuNpa/QnztXpv2+SpPLoxlXBZPCYIwdYD0OEBZISwGxtm
RW6BQiMsZ7wzZZkCu4KvZgBtICgC96ZBcWkUnIBPsnnOprYHvAewSZYEW6zX6X6xDtKAyhC/begE
8pYO+Wi1loaQXdN0InSVmwl2Qlj/q1e/PMHTw8LJIkwbbGhCEE1G4uZ3PFuQjZc8uTbIwtTPegGK
VtZvxwqzsjNCgqa4ucyBUngVGpu7+lgHskQLKtQaUZl5gCwey07KAsqNTYUaPe37tbcW8B5X3cwU
sof/DVpCIAabD9jUdRq73uSxdSuOPtTy4kjlKCK2+ljJGCmerMETXpsUniPbRhissKK2GRgkFsgd
tfR0mWqbbO9zp40SixYi7JuVOIaisVXldThawv0I+37hBDK/v+fyZrdWZOLTwiEXPJ5heE9oR36F
5zMFJIRbH+VX7bMC+myif18HYdxX+yexTU3DK5fTl2w/XaQONVM6HOvYPqSPSM6er7+zChJw9OEY
54wGtTqEwcURXmciIEhYJLh2jw+eyx6fNSrlFRPYdX8CCbxO7LFdrB+CuHBW2+JNTNn33iW/7sLg
yZ3opNiDQ6jWmg/soIt5Q/PyJAfWYF/YMoFD2kUyF8SsuGvPA9ye2txA5SAbZRZAO916J23oATWf
Iqm6nhsUm+Z36ZCNxtMLohJW7IkCDCkl+PQrCse2NNrNAiOnCG2YsEcCC0+oF+e8RAZc5Ao8OvWy
PqpfN8lymLlsSxqCf6hUbSEyUeqz3DNG2aT6osxEfjRMkin/nZaS/Umbf8IgMs3FcWR/Iih+4eag
ehM87CP91FItT+tSHy8a/llFry2Bhc6nfeCVixxzkwVZpQr+h3LXHra1veypARhNUjqPQIDDv0O2
RvoXug3gMC9k3/AezQ/1tk10UEktuqhbkR295mNaHGK9tXMyL6dyqLyoapj2nwyftnFASS41DMfx
NrfyvQcM67wc79z/pfOQ4OA0+zp5deRkuwwXSZmdCVHLc8HCDtO7R/anovvZWLPl4DLMJS/NRS5l
kgPbr7CKGN5sFLdhLE8XWnNDjxLawQR1BIrqHiIwI16OPMXGuDPbvAhdDlZ/II9PcEX1Imh3MAMw
T7f++MRY/HdXke7xDOXaV83+AajFP8xbXPHJOkRJW+nApjpjF9egHH28rmjSPV+agBu9PKooGIfQ
RYL3nseM4EgNO4I19GE9hkxi7QQPyepsUrUyNcM0f8gM3fFkoghZmi+/uBFNIDMqAKToMjDTZt3A
p5v0AcqMDVYjqSG9SrfG+l6QPXlKO/JyeXaFT5tH3GyGIBkMi9wbS1SdRkTqtx9k16y0Ly4EMI0j
mJCjms4E3n/HktyDlsQzuHwCasIWwn+v+3Cyw7VNNd59mFMYZWUdgeF13clS3/MJQHqbuKeA1I23
b3X8ZiLSXyBFB5b0slVcYU/dKI+MKIvRgbTU+e54PYEFkRWcHTFSvDHewtqkIK50ye5j3JdL5vtY
g3s86dvsgxO67nQ3okadtYJeTEJnbiQa5rCe4RRMSJfmblrxEOOOE6JA/e6cqZit62OLR3R+p8R8
qQRkVp2Eywxu1uc/RAo7LKN5ce7+h8DZuQCozlEjKLGCmSjfOsjH56z5t8agpjX+Pu8BozVknBEB
7UWjtNktqpkEpf5uDjNLWKograyytetOdPPX+kyGPFF7yP2/MAvjNF3XvPetct27XmUkq48S6XDu
lFxfJpyF9iIl3+P+0/rZhPjuaB4qYYaFovQS2kVKrDcTWzMpYOxR7ssw04hHXbLB5nbKE6nJO1Jz
GqMSRn7tr2VxyoRx3wnDpPDpCX6qurr4+TzGfx/jhe2QTvwo3oDP18DF8vhWB2hJFgctc1s+Y6ru
NdhAbL7zsuHpeHHGPGkA1BEnSONCQqG9xtQ8mWvPUY2PuJ2uQbEPDoMq4X/lm3cEOf0RHsR/TjMM
4oJZus+ybsf1jVYnAazf0RTfMKrm6HV4fQurIIrKJiqS0nvHT4j3LiKCuYrDKT1wz6SeEM2qn+DQ
0Tua8LvZ7vrROHYKzFUK5Vkd8dz9mzqcwiYs1fEQY8SGAfdD/BTbxni71+TdIoXwpvz/lzqyJGFt
rdyKdWIJip/YB9Ox8KYSqWQzPPGEydLSvkbusqf0DdTBTbX3zSRRwTWh0aFZcASp+czZFg+doE23
WNVXADnfopOiXe6J2fB5wWwCtFliGCRgQZ9VjFTWJneDZVmlmCkTgO6AgNyUygucMunYasyQDa7C
iiOzm2N6EP3vdE5kLj1IcfJ5XD1EO0Gtz05oX5tDyLtHrO3mlGBk+M5hNZxpA6CkSjhvJlAqGr4K
nt4jFBpter01lv5sEoR8zTUmd7mfAlUd8Lgq6SqSEH0xoIO5m3eybeh5mDXi2Gzdi82OJ3/cPL4z
8VQt5e2z3NoGJwXepw60MlD2tSH6xWfW9qNNvUKFmLULRAQGbGtTwefAvt0A9fbRxxAB/zFiz0Qt
/wDfz8qeoAgbSTy2GcVqy6u96ian8Vp2SLopFVbG9dGY08l4xshhtqC1k+XTfL7j86/LiAsQkGYn
zYBf+ZrW/mMgSCTvlb6lqHEDzPdqSjK/+oFJZb9tOimH+n5VUIY+3QHRKooj3PsD+KjJahHKART4
lbJBuQo4F1qlYPhZrdDbbLrrlyrxUlBP+fAgn88jd6D4vD0ZPv09kyflnycLrCuJ0RKkPmZtgQKN
xvP+i3b+Kk/ZJfkGhy8Gx/uTVMMvFSQSRad/Hj4ujUPNqSFBuQn0ote8yFZ2Z2n+vqZlGxxdbtW0
/OX6up3H//za+kjkE7dfrb8dz+kPXg0hMySuE8iwLVHBlWPqR08CfgOFuGoCYGlZnYT4jisaqFiA
Jx1wbRAP8VC0ECaQq8D9gobRv9Ri15fLVR9M9LWryFRyEuQc5sY4fvUcIVpeZl+Wil4z9wmIipAc
bpFTpeHTsJetuesxxxFD3SlrUA+Nu6KdHxadVIVVK8M/D3qKRqBDFHwoAOjX7Kdjgkwg4hVnDZoO
phRfnka+G01MG8r33t/HE4BvdlFycUyuhlaqFWJYf6NVa4uXuDi5Lm1J/RehlUoXhl1YzuXFKeMa
ECc3JDnQqKQB0qLju/BdcLxGamF8uRw4GERInhE5Y3f0DkA93r2hCKM+dyURYN0fD6wyzdZHSwxi
wpevWdgcGnvICt6uEMfjllr/eLykSqpBifNUFke7N7IEow6Bi25uHApytmuJ487cxaFzmrxY9QYG
S6oeF4rae/pyn9m7m5g59XU93SiPAOA0ZhTP36CsCjWUar9mN3LEKTsXdQi1e6c1LhRa+zbjL00P
mqtKap5lyqM31qC1zCs9vqjmleY+EhT1Q4NzKvdeqKYYTX0bIjlzGwn4rYEkIB2HmT4GC8qx9iDG
Lyvenu/4oR90M470bsIzklpSWZI3iWNJPY2qsaaKc/u6hudvC6RO5zjv8WwvwsNscwOI1ZIfTlBg
P7TYbKjGXsSzo27snViMojHnP72HhN8WaukCL5vblfsEReW9Z8Ypyg1crPOQpAiFGugzT5Da07Jh
XdGeNsH2AR1dRoX59kOeKCO0GSzK+SgNnIKiGh6dOS+tc4En3tvho5xxsW3SsUTerpt2RBX5i0aN
gW27OuB8XyvCWDEus8HJLCWkQ1aIU/IkEtA+mVDEsh28i37dkqhrGpuKXmvggH3Wwa/unlRT0bRZ
94BQrFiiRqahb9AE44xdpSUhFMRCMare4riizEwLLStzYx5RJJVXlqr8tODWWYqL4goBN//Zrfxd
t/UrA5se19t3hfmJ5oNstNL+ESulsxN18pR/pv8Bt+oh8BpafsAtoq22kuCtrv8ZtfYJJUQ7OwPy
ocRvwc3c8MI/aHcAsdhMkcPyyQVUiu+Xg7jQaWbMVwKGjzWu9fLmE7j1c+ZwVuzIqcQz1jhXb9mt
yIEo66KEjuDytMpXSPsAqeBRdhLRGRhLvYpwk5h5GI3qSiq0d/pPOiEQXl3CaNebeacnrXfn5In8
p2Pmq7jbREe+m2f9YeoDTS7m0TK9JA2g1KzWDkXBY1K2m7wHSfEJt1iNAMpSHM5Qp1zxUPikb057
Wjz+wbUMLDNir/xm21A2Mly2juaOFKzoYgEjByxhtWYOEc9tPBWzxhLhTP9eOrDuqqPYUnqHp4ak
jOJaKr2rep021ZiCCKdsDjnqQ6rXWN6aKq44RWUvGU2qUDjjUIgSG8hE0k5ZqF0G8C21ynXiJhZ+
ZVJjr0elNjKx2DgnmfPmR+GQTHzjhO+9aLnxd3wWR8ZG4WjlgpoChvRezcGDVV+BJQnM/9XZcSss
miRliw+32KHXHcYzaWMa07B/0+Shruf33bFzdJAHDbotxh2rEJUUr+qN5nM0AcYvC1F5hXEJj8TU
RcBzp/dWjc4D8u5U680b25G5LvdddcD91mPv9kNVRCOjosMllg0LrTL5mDC37AQQmKfw4gDYS8kV
5LCj99G8vhOx0thm1M/3K5/RtNFQBykooy3HR9LpyGFUECENgM2nh1fqErgtAHdNMmRnjOCkMGdd
G5PWrYnAY8QZDhBH+CqewptWdYc+zH8dKu6NTZIAqa7J4BUInuafbs71gEtnFbrNzw6/4VjiQgxl
6mzrgZ7PGjrhLtn59DZgD2Oeby7bvcCa6xklbwsCf/Ve3UFU/aiYsxrVoVbu83I/vQ0vHjU19snu
MdJu3EhmOjc+2TD2WlKFLDMVqdylW9TTSpLm/o48XqNLQyWuln6BgRe4XFKviM1wr+JVztw1Mk/x
xb7Qh2JoUXOGj2iqVW3ik7FG2m/HqEqHllG/gt6gnDPSPXHl/c1Z0bUpJ4r8Pf4kQf5uRJj/nQJq
4/PLaApOvmKpoi180VwdT9S2aRLndeOjLCtZ4ns0u0g5CqveMQiWjUIQRRWgCJ6XsrOX7RAGdE1f
sxDYofr4egWfyI9STir0y0B7ZD17UHkZCK0GMrn/InNmIs21YtoECArJ9t/LzWP0hlBnLOyVBt9O
G33XIotQ+4fZoLuFrPerrqxES965P69IxmX+TZiU6XY2kk5Aksz/YwPF5e+NvT6zO+FsfGHo1rmk
RSTEIOg88y5RfrBXTmXNXRw3SKNlzxmqD6URaEjC+YDTDob7ZcyBBRe8iCfGij8lP6xPaCiCLmcx
HXIbXM30MfDE3GAFaH6b8gxlkNUYDnEgsekEQcn67z5FbTBicCE1f0PiT876JA8IWI3nQM9s7iEM
JeySBIVPeYXfosgqGTK7LuIm1wquKvcr2lJMoHESTh8FWte7N/fCarfYQoz0knUML9XZfBYCaoIG
PlMQsfNZENl90w2q2FESWmyyqTIWLfd1T0F+Rb7KUg/biIui8PTkep7wbxrdgAfiwWLxpgWFxb6u
JnxGMBf4Vgo9Ey/zZ/e9aS5jWAfcjupAs9hua08rqe+g46x2uR6Y7mljrXat7ZMik5fge8le+bX6
MJRGqn0AKrhyqpuQLVyaJkKBTXhWKiLHj1vIdR3k3NgSXc70JeZOsc4xmw5R0ZEvN9qyeA0lFcna
w2vCPAClcssAZ4fhvZ029ipIi0g2bPhMiJ4U15kR9Xc4So3E2GoE0/UbjXM2rOPYU5QoY8KJxRhx
w3iuxNDp5ZMxtfLod+xSGoEO15hSmfyS3VYcHBWNS/CMQJXUo/XHSDl7AWP3iMStPkQm07/o5dly
cuc5AEfsmfE1Yo4/M47CVuBgjC13wfMzrVl1YO++OK9teqNjd+UxvQM+91kN6w9Z9aKT54zWCa/L
6qoBw8015WGSykCMGtriOjCF1H44snJUjAUjB4ylmvgNLrbS0dbLIEqlDjwTundR6V2fonRQPrRS
YV3nujlUhfa4ZEJr2bLQbYZ1Vev7q+aPQlOxDCu1dMNCS0hdyEB+LN6x4w34LqP0M7zPrrXx+WyI
HwNFC85drjLBjb9fJwgxuH/nSA7qyjHZ3ISdeHr4SBcByaD3QR/wAcPdUtA6qJ5f+k1Yk/KxRaBy
RRqoaKjtKxOjK02rBw6iDEhs2/RMH6bVHNVobDUZ/WadTVj6MVS97KWXWaNBcAOhCxHGt/NRbDI2
BPFYBQWovEjCIiHoJAB7651X7Mp+++lbIVP0W2VLGB6d0AhLD+sk2dqC2/wtGoFymUqWmpE2UmT9
KKqbsybVlzW/va+pbMQSaj/3GiEI2M2LJDquvDmKvg+WJPo5FSrVUwGrxRa78KPURFA23mC8NZRd
FF9uH1tgxKTYkCNnKsS9TNufiCDsJejZScQ4Gt8YxOcqWr7LWeOziAz4NAKNiEjZqUYTBtibT3tU
uy5aGJvDFD8Wzo7+Nj4Bopt9KUqYTOaX/MvnBH3vs/QPeEwwBhK66urVRQicumho5O1AMvSLv8gs
dUjGnDAe0wUm9StNALA2lU1DfQ/PxrV2Mv5ydHZy2s7TdSV1jsYgk+IRmgQn5iw3euYcT4ls8OFQ
mswGEky1Zdpc6ARioKCE1l9/917HxgOFFomyF0U+MOyjmCR4+7aALYsC4jBt/WAumGPZ9mwLBinX
2So4/ZBnnAqMxZMnp37wQP0kwaIwvUch/9CUZ8KnuB3vY8UmGgJo4NIs0v6UpnnM14OA+v917j4V
vi1+UkKksj3Q+Hh9Gf6uR1fej0CBL5bfx6HOJO+Z3I6C5SRyhz1F8qqFxdOcGet1y7Esvd49bqrp
ocHr5Is2oIYAHbInA+MjcJAF7wSdhNiwZYyHdRPVYpwc+7KAdO5pGS790kpoEwZ/Y8gvFpHEdOKH
+q0SVbAJuOvFmcLS3bB6aiMMyCkB9ueket3QYNFOGs4i/MBP1zsH+JODF3YLWc7SHIozPY8eJH1W
UU5nTP2TWMcjtl0rKMecMwrO/TUqlfgZiNbkIphfo0s5UW2UU7PBkAHOYN8U4XkLg9IjgkZIDye0
AaL+R27Dofa7gayIxzyVw3E4Am3snlFZ6qxxV+2VDUwLaTgwHph/SdMf5ILFdgcySxhdogDoay8z
fDIt844I2qX0u8VmmfIrpR8BrLVPVMTFrv2q+zTFQ3c1A2UbDbr7MFj0Pu7nWAn11daB1lDzfgHS
ARkArPckXtNrk964o+z0LfSp+C9if4sJ+5rmenfbrDUcdVOUlF6fqkkz5BTgHx76/UTQ6X6jpuEV
Q+gAHyJZu5Q2l6eykXMMZ51cOqJSHSuJqrKGgqzdwx4K3JScQLin4F56D+fXzfQeGSW1/txCNreD
kM8bsXu+yPz74MFNw1XjuptrUrffBPS7jgCj4MiYeqg/T9FqcSjo3PgJky3xXebKRVLrtjc8zOmz
AJ/w02j8qRvPPN0OKKWN7P2f6Q6hvaR8KhyC1SC63WB/bbVLXt0jlw77c16ta+QEosOotPO9W87X
kGg5HQrMIPr+WSRjqykIiwxiAvXSfW8RDAwakyEMw+KnkPVxT1Iev/sZ8+iR2CrpMQyw2GoUgxfI
YYnd98NJzwx3buT5iocXi7U7K83Ue/beKi30T3JWqbOLAlgwIVLV2UfDFmA+y+QDCyOKiIGX2xA/
D0+EIXkHhSzOlj0B2uA45pyJ3ghnd/QeeV6H1wqoR65Hd/FruoX3wEUw3TTnDiTYYfllsgqsGnkt
65BpbREoAnN2vzu3dBH/laccEIuM56H1DKd6DFRlxX+IoY0RpPx0f7SgpVD3DVcKXh+NM7pQdaNh
XgYKRlJ1u1z6Un9EtK9SBRtAAd9Zii3dxDbA1obYCkgQ2iyEjsdMspd4iuSiZJkJ0SxkajgFFhCI
GvcF+KcSObDIuLlOMe2PLkYfUWVXtfllURpDYaT3OX2xHdnFIEyhSwvZaypIsawiaJLJVWm4NElb
YDg/afV7urNkXOF+d90uMHQtJp6QumPw46hRJaG12kcrNfcsYLsCGHdv1VjED0TMt8j8q9aIcd1s
nVCXvMytIDLjWQjD46hqz6pbULlG300Jp5fOstROYeq/Cr8nLchLOap02nlOEdaWuEifP4SQTRLM
vezv+GHa0w4cKMA09xUHuaoNMf2xqJr4iDkm90IhmsZy8a9KmBW6yuATSlHmRNg8U/bnDJKKTA4y
l2+74IM9TgZtrqgyxj1Zxk70KIC25VVbqHPOewaRLsD08Ol+Lik4NpUzmhWYEpEJGpJH0X523mrz
2flD0pk1sAugHzAChD6o6JrrAKPl366CclUF8T5nFskjqjwyMcdsaLTatfUsk+dEgQm6/DKXhKoX
hNk3A8iMsK6AN1nxc5EToPD4Nyam6Z/p2JZ7MagYcdxQ5KuKWuypvEX7A934I6fTJb2useVqu36o
tFDjefiL6e2leu2bYDh6D/IdjWo3vy+xfeilgWlmSwTrYgBY17fJQrFrxvkcZxjbPzUotHQB/q8P
jaEvz+4mvrK6vWkWdjKB6FG8zA1EabjZtRtOaSIaaIMnhyJ5XS/eHzJrAN1m2aJbS3CsxMmS5wi4
fiM1Qn0ccSlr8sDkCIPDb6diWtMwcGCt/8N0RNDeieUKlFHx4jYpS1KKbWONxfVteJ6w6NBL7+0/
hH41dt2dYtb6SDJzXIssYcym74Ybh1vmkCTekbMJk7GSBfAKqAsnrxeUapUFnLsewMLvjkU35zPU
Pqjra2uPEiq8hssqSVo2GuFxPciRnhtty7YlIeU55CvReESPpo7qF7qmOnHz72c7rJdnfNs7WTzp
f17opPRqW7275xa2ELWz+Tt/GW/5kHkuvG0TwTFHbEWQ6W0du32PKRHL4AuAKIpbM7EWINitGPoI
mV6iMPKV7elrAmkXn91g/KyG0CKNdJuGDkgomPjmUo5da/bw8xUK0LjYgF2R+dL0oRl+NKrZoDl0
wtVSL4dcwJi0ampDURDIeZnRCjtFDIj2x0a0kbKsNQD0ZH2S5TwOFx1ArZR+H/zoPXhymyXYGHB5
px8tM9DzhA8UkbwZmTIFG906+XwURhi1jnRa2YBTGx4/b/uMdghMG+L8/RaSFfn8smSuSY/UMOJB
Gd+Pf0phMq10f7kJIpKTdXCCNIWMKKH4KzHGojFMo+KRPwwcNt0vqH+vlOhgrrGhE6FuuamzoWfi
jFj+5YLNUMVX9EmTCsaAaBfZ5MbH4LDiEHKho39I6DX1axZ3d0dwaAggy4YYpwM060hXkTXd42FZ
zswczWggSZkBCMfg10XJa4CSklN63YNALrmem3B4z8568qdj39s65V6dZ1fvQBj+DDpT5ijTSTsO
wRAgbENZPimNXAYKUAjAt2AmO3Shx3KXUCzb0BMfVyOMse6IlEgjK2JQxWeZKSlyfl7kbEwJuVBr
HZIFSIrbdwV3rcNgv22myglrxkDAng1Ydv9shaQYl7ulSc442WVuX3wR1NxNJpvcT6xxef6ykq2H
THNphsVlYI31ftBqWM334NyuA2F3dWF9tITV/dH9kgi2YP2c3H4VXyEV/a4Ke+Ous1k2Qmxn7hhc
IA2QfVQaTpEQJQrwcNDC5dtRIDSXznyx8KaqDoDrOuq7xITOHibNFOaj+T/mzzHP3px7jFuo3oLk
24yAASkF3eBIBOgT1mas8BEx0qsWflNTSLrzBYZxcZZsfO0kPC52p9jt0fwTFUPaBA4AKAg/Eqoe
6z/tm3huPNXjRNRE21D4uOIeDVN2cYgVSNovqj522SXNsTDxN4XzJoRC0TUmRt4LZC+ORd3F/5FJ
YhbNSMsVnQPlWqI8bsPhNT0AHwnWqvG5jQGYM/kIt3z0pwIo0Q/dnfouAF//2SMRhmcU5dkrFQrW
NRgevSqctFtxV0FbhAVRKNnJeqHL6kngtc1uwTFjtKakbkNklfpk9Q7ZpFR9p4Ut7TO/lYHBrrSP
Q5QPGIDoGYM67dBdaGEoQXrMLw/eOwb7uuXzNGE0Pvon+HkCT68bAfmO0mMsQDwL08uYCS/ar8Fm
qMAsvAIC+lS+qm2LkKbUIqWKuac08rWTv3ZtWjQzrL/E91daOXBOCBx3EhJ9uHIR0fkwAhIyVZET
74yA8DyaUB8hMsmhzMOQSBcUYRH//xSN8/iEF6LkBin4Fv8jlgVE++L+yOx12rMat7Fv9OdfncF8
lfgSTLe+AsoI61ySL/X4RMTnTzY8EEkNKwaPiwO/Nj+bpZFx6OE343MfOfFbDmZXOq+w8YOb/eup
s+k/w/wpDqR9X5dvyHlyesgVuZLcJD4ei18XTrYG89EUwFjcGS3Ra//DcP4rNlqrby7SrYRPAh0K
ZQl4MYDXY5GU2LUgr9ddN8i4pNoAW1u20gGQ0/VQPVbFz04TU8pFztJE1O+RKNw2WTIVybDsfkxu
hEUzOHvwm77cvgG1AKhGkknLsvdpZe1QacaYPQ1fUtAhYVIej67sO+GVkLOybhfyQqcsAxjCOImL
aNyQKd/VClsBd9VdhHizrmB3qni+coS43/X8CoG+c3dN8OYMk03fjQMFTaXpHu/XXHTJMLHI2SUr
ueErEuK29hrrV80KNaqSekytvrCpGjP6bWw2I4iWIRwGDuoUviHj5PTuep+Z6y8kp3mx1PkAmkkt
BLpE7As5x3OztzochDwhjQDvzmCRNz/5jMIJPohBGeCkxRtk2MhtaFcCq5kvBMuMte1y8G7ulFgu
rQO10pIp8jxIICFiMMkSB9onIdX98PMbFPrHbgESrpcOewznw8toHL9YiVt5PHH5XISAUkANMreC
xtuU9ez6Ua2Ibh1cmkbyUzP1UDLsDUErhugsuhKKPUVRXka2fMJgP4/m9N/Bwf4l7w/xyVNxlzoU
gEkpYkPcQvjRM77foiB2KOyRiR5G6pAdgQTxXYvIauocWbZpRHTjkFxVJmnQP/JKd/Vli155QjY1
K8+PmP58ycF/3QEsadmKWL2lR+qDlIhcOvYA8j6p+UMS0/I5uOuIm1DyrStWSRsYzKGtMRkNJNSE
NZMvJiGZTq9K30g+HIOIfnSrXHxCVZ/ovt0EeopuOdnsg8i5V0Re1+N/RdsJgx6S1f6CbzDV+voO
EJRXL/pL4F2dEvJM9ese4j8YhIzaW0mvSAM553BeNkhDkfQ3CprdulysZyNWNNubliZ464KZcNi6
LtVnLUcXbQrVNh4F1GJ2h8DGQ2qaHJorQ7D16/ph2mm32r4OU03OEtFn03LTxwOvUM4yH3+ToZ+1
jdP+kwi/pnjBjyqxGxjQdKz2S01FQqqVwxxx0RomPBAHsH6HTKlWiMPfXSswlwrymYePiLRF96kL
85F81udtBzdBG72ey4A3sGn79erGwKYQZKJ/9yIdpUxRjcd9PyS4Dyv7lDm780iUWnehsPR5liIP
0gHake8SbdPoAAU3SHogQGcLH3EzGLqcZtLCe+26443J9l2kHt0tK6BASlFh+Oc5Yd5x2Ex+oU/w
5gGbIcl2ZPDpB86XeC3pf7QYxo7DTVYtKhiCO5HZEibE0ypA3cMYW3hosPFWi0vTKzmqWFYe4Ok2
pyuyUYZL43Mqe5sWyu4VID0AbscwfAubzjZpu5ApddmjkbTb6h+EZgzmnub1PGQzfY2PPyVneooD
iVi99+tbJUPaBKCDeQYFuHVpsy6nsRtJITrxFJTUbNIhA6x1d7R1RNfHeov6fpPE/9E/VIOKxVoQ
bIDStHVmvNZ2tKGxOD79HP8OukY9BEo9+PVt5JTOOowc8TdHobd6gxr9VpihQJvCiee8Sn5Xfj9R
U7E+W90vkdJwSPcu0w0mTvltNA5d8c5Z3JLqmdTsvODhHUTnXV8YLzMl6edhw+cWFhTLznpTqnFm
KXqas0vH8XOHOJ6Uw7lGjjyd8/JeObIeTu80KkfpCyA072SJMPKeLeqvct7yLx+HYcuKaZae+1qN
AnSxP0w56mDLSQUZ5NGQifpuC13CWreVaO92eQGSWRnhDSysVtwd4ArN4kHAas+3iaq+kEAJ0QoL
IAgUKiawu3UPRArlPhNFU9Arl0M4tZulicEguExoeKJVggHgaiRSxpKN0uAXdnnEDo2nRDaZvpbF
YXhhCyWPeJKtSjoyX14H20BBX6fX2RmF3EafAUFC+eLC59PxTdXFIy5hbRuMztprkrk3BmS5Nulw
PBQFBKfFzsTdKeeSjp0nES4mPwpYjnjQM+YscCBtEqh1qzVo8UUUt2U5+lFerL0N8b2k4L8JL1b4
yDhuTPahWL1B7/K1rhVMen7BI+SDgbXBQIEiXN7mSi09ocxeuTY/6ViYHH1Jgmt9bTFur/uC48ZH
L51nyXb9T4aSRMEcwA46qhNFnP2LTsD1wkQkzuwHAc5lkG9W7ZHs/NuufwwUaRGjPjvwGhADtmYn
8ye0EalnjXLBlMaWwRtTLEKIapa1FceAO2Fc7DXdDdDM01z6fT/g+lwzIiwzjBEBcp34uDV8QiUj
48UaIFw7HmwrxQ009cZ5chPwVbqJSMEFZAJagNfeziRl06zYNFYIb3IlpHnk9NAsZ+Kbe5iiN6Bz
3d/CSamsBYR55pjRmFnptOZ/GTR0OIOvCrPACiInc3Cn/GTrZustVpcXlL7uvAIHNbTAr/y7+7Yg
q+7RiZvzX8YLi4tXq8iKoX9gxGktUxRXFQJEwA6upwGSJbq1fFiClh0S0WHam/eifVUjVi2vrSB2
w335JoAzmEKPNbU1VpdslT+XUp52PtNUqrYdEADYEHQtCj1y7Dy2ZScYNjdzX+JBqAJTD62KM7OB
jzX+2kNt1dGGLirQDqcMPcWI0yOblSr/U4fKh6Cd9JtqECQk4tGnxyjLkz/9aOz3HXsbz+JE6pqU
+a0Xw8aVkAmYIgjMzkVwCh4Ea354aYl5HgEJQxH81K/WrYjxQkTKGlAKOatFJONGDSSDxipe8niv
lfnwrWkZxRL+AO4HanbZiaFcdwF80mEv2BjBnNOB6fZco8YiiO8bhiEkjebDi+17hNMl9mCqzSo1
H1F44dGiGX6ihTWJ1CdF9LwNIVx9Ml8Knk4ETGvF6mB9umVdf8E63D50nqU79LLsHJdIAuWK0O3J
H45Jkm5DtbNaLbBp97ISfAls06eLe4FqAdaXOZyk9TVlkYyd0CcwR0URFZvg6yPbGzdZ1YLe5Z4l
AUgsSXAc7HxY3YEKwwkabYvP9LmFPDY/zeFfe8V+tZQ/lfXp99maH8HN/I9rLFJRcfYf8w6kXGcv
X7qXVr2nonpNPcldjRlXn5l5xCe0aIOL316vQrKN68pgFWVmsAskvh1fyz+/8UbaMXItKg9QX5xD
0MfCsfsWD34ymWUnHOmZuB4OXQPbiq8ej9Dpe0p7aIjaxaNJf/pmC7mbuPYRlvomMBbpNLFLz3OO
gMaJIy+Fc2HdmY814g4441WzIhh2NM3+UFClYNqG3pa6zmoUHFODVxIcOAQMKMNKIYc99eD2n4aP
n2Et88QcAbKjJx0n6WT0l+cyYbim0m3hlA+5+y9lIVMCpzJCPt8/LB+bbxAHnx9LbSE/wfoDpGsT
Z8uRI4qefmZckvNBL+R1UeqUkM2dpKYOI76EsC2mfq8ghdMEQK0pgwqyNPdS97GPZfSPKaRIpcbj
xoWACJaXSDXU4Rt1luzmMYj5M4Waof+YMLqzb8/1dNJ9XHjvGC1pbiySDjZF3BBvOz6GR/i9WyjW
Kz5YD/X5EPwWhUbe9CxdR6B9Y54NwXaRgap1PwqADTBEktAodgzYZ9hlmVmSw/+x7OBVvc0ZxzLH
FQrQ0MmhU8JBIFmTfQPmkMp/aYB3zajnFwH7Z6eGfBAqKlEfr/v8yXP9AQ2HRakHZA2AnyAMrWmc
DPnaUpevd+SXbgQPycR/PjEnzkio0Md/0a7Sz1AJTBaLk23CblWBxFHHowECSQU7QPvnwCtyFXew
JvjcKrQunKOl375zOLrmxT1HifnC2JGaQhHy7A3GDRf8D5mP7FxUDMPT8JGyVIXBmdZgJG0mthxo
VE8FJahwjKFdQyxlhyhmRZXef0/ydTFVzSW8BJOBCZVH47A7/bnf0+ymrzyUP6p8rF70DkhaW1V8
6Nz6yWC2yphUvUpCP6DeSHFgGH+7KJ0A85W+TpTyrkJLHzU+0t33IAeVZfwJ/UfMRE9aZKUFUL8z
S9EGOaY+ygjyJlLokgkPHPILqwLGy0dVW1RN1+muTwUp+EpuZXbt1KyS/Krb71jeF+4Gd6xDS3Q8
alGQ+A/9whFeKD7qpYpiIHMUgYTX8fujo9emePKsFXprBXiMfYTq7qfkzvPJnBb/8dmcP/6QI1Il
wuy0wOaWfWAWY6zT3ELisM43mDLjKjbCZZPxn+Dh8Q+URD1aSkprwf2PiQn6SicrHjyk6yTwoavs
9J3Ktu3JqrXwIgC0EMGwjqRbHFoZ9/qIcyaWsJkCNqgsbvMEIKwNs3phWxe9uXdRCIvDIf7WnqH5
jN5lhgwbTAdmkxTyMBqHdZIk41DWloncSRQfktC4sgTV1KcieSor/PctQpCvbiHFJkg1jH6Ywm+Z
+r907Wy+so2MIkzyiRNyUBwji4SvXwjmWzPOCCYiDtsUrq5Q9BsyL8+ftvLQHEC4FntHbb7DjBWh
xjB08+dP6Q5Ab7f/GWvO7xQtGcXRHXiWMpoxBJcyfwKoDc27Tgi83wuo0LOvkRjkkUrZMXFFoQ/v
oshuwf7o6Tq6Vqolyr4JR3zkPl6zpw7JNp76SUT/o9HBE3zjEXSQv93sNdiQ6NtUqMyXe+7/jxmg
pX5mMN2c+QqxTPKjTENK7D/WePVfs5dR5Xz+2YvPk8zWuV1AHGx+lw4QmOhgP0BwB+/DIDZ5WhTh
76yerAIvl568SmwqbIGu6uWFX/TMw/evRliFc7Qda4umc6ALcTIgWpY/nweZDUENbs15rGMUvRCA
IVia/geozs+HOjJLhUslycJtA0OuhCfi2Gj9uQmG64f7AjDn9g4+PBU+zMieYdj70YmJYXogHjRX
m2tDGrmZL5mYMW1O+dNlwvOqwnfi18lRVDSMS6tjeT10ZNxu4e7EanYZ8im4nlVWISXg38A9DqEg
IT4LNZKSrSNiPUEYTk8K8+kv/J0SOYq3HhY+2nXP9/6vuZ8v9+aTDvDwPyubSJ0GWaReWMzg50Um
HBqokCPYN8AGL3Mt9pLNbVL/9Hsy98zsyUpvpiOvEKI2sH7s8K35TJQLWy/gUgEsEEkcbGsx+X1d
PoZO8cODTIavaMhLTKBXAjdsvC4JjFPeu7cV2croh31Xi8Uj2l8UGxEwCofoGAtycapz9c0iJBQV
WKnuui2mKb45Wart+UtneXLv6guAt6UySyyT8DstFEvT/HYnwLRVJ7J0MzCjYgze22Mntc4TDWm/
vw/7SzyOoYbftOtvF0r9Hduw/EJ642E4gi8w4j9TpyhZw36ul6S6Hf7Hr/zgp6MQYIncMRm2Ivkc
fdQYCaA0MwWZUtCwjli4p9JTd7qXps+arYgscShQTXSqNDbXlrDexDldVDtmQ01GjmHZdENDUT/B
RnKvFM732QWINdV7aUCqFlyJ7PBb7UVI0hj6KA/bndDr4CRdTMyj40HuCkp0wCmwgoa89+oVeIV6
v+wRdxLkwDom3KPJeO44zb+Ex9gZOmXEX5HeodWOmIJ+xEMJwU6jB6GKmCoanYo47t1hDuXwPynE
weRyTUAKVsYVaMSo4ye8xJvX3OqmvEcvgPFx5bKtDSLghPbM6aH+3t0AOfifHk0ZCL0ZHMASYrao
i+trgbq+30UTO3Ecdu5lJj5EPWd1sTv8qVvRYqH9bD9OHr4LmWq4go/19mHsuxzNX+GbPvRSOnmP
eNDok4nRgBkZhLgDx/QR44aANBw7L36KDctaYddlJKGEJxRrY1zFoaiY+hvkclVPzJT8zecQhW7B
HHA/fXNC85FMbNr5Ovpo3JXSKCN1o65SW+0OxxEz8mJ7bt+YsGfYmy6ornEMmZBAtqTgpymGH0Lz
3LPvnQdjE+ELMkv9VNmGAYrxG5u0GS3+nwyUtrOrAexv9GTFSQS9IT3CndE7lf52Lpdrcak8JZkc
5/L3TKNy7PPLDUSkUGSa6H1pkHn/kjQjpe0BhQSQI2Jo3buzNUxpOrrYeR+bj4hrrkbyDl22UBoX
/waA4qLAUP0MICVwtSGt7/k1sGac/ts4jrSGaAYzhsaApx7ok6ZkCeEtYPkDDp1jAyAU4KyID6gJ
c8oGIK0dkZlZe7WQOOC1WRqFpx19hlNrbprAwJHZdyutBgwxXgHfhm15FbKDmXo+Er//r9oh6og0
Zd1uGDtbgkXw+A4YunKWXCKJtc57Tv7dbqnWNgMOkayYUNUzk9zEtqG4fLlh+b6LQGTc+lZabL4x
PHY3o3uimr0CpASPxupsN+rSOr8x3y92+SPbEzQ3a2B6izOx5irDxSRVQ/r6BPUk0tqgDt8ZwE83
/WBBTFqACml59cAgng08dvYa3p+q48evgEasnfJEG4IpZgPT9aN2Oap0tamNxEblr15YbRbFzEAr
LwJarLJANjuRCqP/aK4n+AcuTGCdi03pBLbTAwlAe9D1K/ushRwVBu35R2fJ0qKlcRWMzdc1Bv/E
rQiQzcas9+oB523gzEpg/sNA+ZNrh4qOPZYP0SQ3uWinRJKyIgrylUNIBR4DkAGrcUQgtEHfiOye
1kU/aJ5ONuSazAIC4zUD9fR3qYGwNxtxmA4KA3hhQtPUJBJxUbUvzlrPVw6gZBrHhvIAyXeQq/AS
qOu5IX4Y1y9hWpkhBR4znFpSOsR7hIlrCGSd5s3cATZzcSq7cJ11/3oSGoY43yb+ryO4pamTxMyU
utRYdPcZR+BnDaJAPcOho6VN2evhwmbqRF6y9OBqr+xhLm6G+coDfSavK0p4u5xXKTPHLRLWiftY
ZGvmOiU2mF/HT3d5j0K4dB2cHVzDAOskJAQ5oW5Xm62YUCT9cip1QXXlj/brz5UUsUobXdnGmKZ3
a3mkvhCbjgybQ2y+HLVJrvlXtqBTGBg6cWGx2HovlQqbMSTNzNPg1l40x8RRsfAzHy2cQBTsbQVl
FFbHyhZVGHXWhYjQlVxFCp5lySZAT54J5X+pW4HaHYZettcSK2+J5IXMvbJG+q8XqWlPWnYycZcJ
umr6E7UzCVuEYvMzXOwM8FDXHL9DFXsDNxl2xHHrTvJ62MT5q1gdycyQui561IN5ZJoRxinPjAEb
igDEl7rD5UasJdUww0awbmpXauk2x6VLa3GKLz6QuzoLnACvDaenpLERR3EqZzdWhahhOpFxsI4W
rJYVjUwvPN/XT/k8RQ2vWsvPI39o4xcH/0d58+2zBMkSySZfuBl3LtEnk30tJvQFGR/Et5TwP+Oo
hq8JxSXpFTkf3vjJhlPkZOh7xayQ+6OSaS6Lfs6FxTGrjBfXPFn/DAgQ+LGDdI0ILxppGaFuAdb/
YW8BbGvXuL3RrqVpOZQTLCm2w6dc0jRYk7gGv8jIOGpjElqxqs0VZ9Md4Gam7ib1cghK4/SzbsQm
PVRzAULfFk6nA8o3tLHi7T73v0OUWN+bJj2NOqnYUDbT81iLzrkVMcZUX1VNcYTdsWYy/E3DU9Vh
hhPo4IOC/30gr1a4kGgNSvSCE3BvzOyT0uoa+nqv41PsUgVpCc2NIM/cR4wsF8/i7kTigstetgvI
iU3nSr4gAfWdKhoyOsHqNuDtXnv+5Ga9ZgsH2lGMHVBnTb6bX/u5OU3UCo8Q6EnoRrLlluqexCpt
QszGfihDmB+wmTnKxYrIf6csYA6h6/gpm6FtbK9PaKGAs8jT8QW3FsBInxA8kHkKiGj4ZY/ObsrT
rc9YpzS+WjGVqMZv6YoblKY1zP7R895wSt8wDnDReAbIjsuU8LFSe6DH2vyUcBaF/6dQFXhcWWQd
HXgvzq0Nn5ORNd1VrPn8sJFhbkmIV9qimnKRWDYCiWNBWqDnoF0n9cbOyMj+IJbmycFORLxlBt/d
1fc5hFfpNbRSipWEEeRN9K93EAEU1IvG8r0L0WhlF53u8w6Hxch9sjrbIVsBu1Via6aRORe+UNwd
UkadJpWTcL41KT+8DvUXJTDkdqkoWMlRMQUuU6wYqNmZ2jmkJxbT/NrmLufND8CE4UV1jZShtUU8
Y/JT1VVB1m/SdAgD2aGwrs6FisfJ7Z0XyGtJ4VskzgXJAHQ6ljeQpmHj37Mmt0Us7cbv0hzw9m73
SBiORuLrYtxM3BTXcqxqxWlHaZKS3YrJpxNl4q+4ObI+DMIC+QvvIBXPzAgp6OVsE9X5b2CPEiU7
4bU37wjmHxtKWEra30AcdMUm4w+jwFIf6jwN82KckmmPbwGZUt9ChOsM3E65zXwt+kbkD4z5qXFr
M0JxGhf+hbgYWaJ+OwxXHa3Qt/5adBTyHtlkgskS7Xh7zLYi2jRkKRMCP0J04quQ4fp1onoZRCoz
cKGPk6rWDAeznUr4IQw1CBetS8IQh+HVY44HybwcPGK6kKmqVAZwVfS1KM9cryAarGP4w+d304lF
UgGIUVP3aCeVvv4CF+J+CZ/MUqGTGe5E8nTdb5uTI3NP/SOhrzk6ixjepBBcJzHoZTIO0hiK1GbY
kLEd7+2NRIK6RnIjI6DIosUYrKO3/7VgzrZB93Mf4BX9FJcvEKbyTxJBw1vkfDUjFiS0AbBzT/dd
kuRhgIZShVS/chEZKEKRMEJj8p/D/+jh37p5SYoiyJAzcYuB1R8FYpIB4+zuwPIpwadHkLACW9w2
9j+mCSOHhbC6Hjdx/LE6/HiZroOpx9AxFGXkf2BV3OEIULdL0S5NIcImnZ44VT8AYjsQZZYk/p2X
VJLZ0eJ40hHl2Sd9kafxwrC49bqFDVO0qt0JpIgydAA6529QEMltgUtmsJ+c/wbi6jnbanyDSFOq
RiitGRumZvJtCfl5bWQ7xm8fRIpJp9mmAjl8DNkEH9GjQX2DJOhn/4K5Xfz1koq3U7o13scTr9JB
jIbYj59aHmUfIZLuFaE3xHHKUEe5Op5smMwEg+3NvDyn5rLfVv5nfRiIMIxvG+X7ZoKoAkXnwAkf
/g/UzVwcghjqWd8BJjvUUAmdiaFep9wp8L1LG9L0KmgYbXSvy/SF23p2xpQNnRHVxfsuvj/tyMQO
veEcC942RNtRxLLbHcvEPxwMa4NZx4EE1p/BPtIZv38Gcobo/jbNnSfKbm9j4z2ql6aqX9fefCMh
Km2yqvpF4hnqPGEoD7lDAI0li31PwMTR96he51BuVpP7NYgLansD7IC9PAUL67jr3yOR4aR0PDTA
kFu3MxP/OYlGryOvbKQzR42Wjxko0UACB0YCIbMqYKSDEKLnLNmQ6cR+EZDQrV5kFSKxxyaeRRaT
yUpjJPQWeKU+p5urihvBoBJ/OIP0w0qm1GgndCbhCU7WZ/wIMsWgcMDPnNFcMtoruvTZVhZYOUsm
C6+iZBRUherUki0Q4pFm55dVY8YmX4XuqFd4vqlzUe1CvYPL48+SeJA92Wr6W1R4c0/oJ+StAaXY
YFqQpr/bYSRgUfaHB/Rl3PLzzw/3jq4mnm35pV+6wtqD9FDzykUVpKkWKyqyojFjA1BShwWnQqQd
OUUl1UHWiSL4J44lOjTHSD2YLwFp8FeTNALsEQjTS9ecByVgUWgSCIadIq3ErAxq5/o0CVApMxFe
XoZ6Yp2BZT0ctIuXnoTWE/pefSOvVCfrRIFqCcmCwylsJqf9RXT3SnBTlHxXnHQX/DQg9iVoFxjX
2IKtiHeSeD2RSIbtQ+z08tOyD9mLcUzorCGMb1GH8wNAvEjxhsUT1/0rmsnlrZxKEjzy1d09kEsa
XxbyW/by2H+eSBruF9owlZZrRReUvra1z8HLRg/euJ06HPfRLpbXXW/L02LOl0VuB1oZoOvrhAOw
qOijYBCbfB6mHg61c3grlV6I4hpmD+DL/9y9l2jzdpnJaR3C1Xijzeu/FQUIUvmCNOQbp23Omy6T
fun5NTC0MvhtCdLkdX2e6wseNxvYFPHJrtwURWK3mXQCk4+vCRwwu5us/eZp6hrxxG/x4sOIgpum
X631l98aWRycIibqJYPTneXflp6Q5EEHD4GaZ1oWEfuYgUZKsu2w1BCSBrnJYgYP3E2CTjldTLMi
/ZMYFVwkU6B+F4VfshJskflkSuvbjBmpTgSsfKoSTUZuf5hfTHbnUNtPMT6Ms6WdhjKO6euhe1Vb
Y/xdmTu0i/6HqtJj+2W36EwNE9aUMgL9b6QWCBEb2JoYgwTjSpb1bDA9H2Y3OycdCtf9zl4+8iyZ
PFqXKnmDy6xOHoY315eaW07pk0SCV21zzK8xxa+U2t/si1dU8+iqkBXv52qRNRZZLXnnUxvM8MYL
7pNzy2jdOuzhgDjBlGXGqJajiGiUIabTpGNtNe9/enkTz5IBomKrA2FgrKGlkNgFP+4ItwEEY4Ah
/ZGR79W3Xlu/KjHiWwxqyw/OF00eXjl/xa34k3Y4qN9yn5brgP3JvrvvzeMyxQMc+CIpRSjVykYv
AEjoZHbIMdkmvOaUbKQxNCeVEePIK9TO8tMx2ZvKbupzEWu3bICa0Tyw9X2++Re1Mb5/ibfxj95u
hTJcEGhp88st/YzpmIhRizJjzx/J4MgILxag+9oB2uYG+H9pzcaGn4pfTmmpM4yBDqnQ3dQLxztx
3mxfc9ueUeL7QfVWVOuQf9YA2BJuOKICOIFY428qejw/fxNkCMea9pAlOI3hw5/t1zBEnbJCPsYW
9NP/iBaDt3LNOvchkPpgPZ5T1sEy0ODIpRN20V6BCMhaQwObS/GzSUxw67N7yMKA2eyiPht4r2cA
dF4RLk1cf0twrINzKFbufMD4X8/GkRF77NhR0L8Z8Of3750ytMpN09oRuZ5UB2vvOXM4Y1wDmelg
huTM6EWA6yH5nZ0R6PH77xWlr4T/XkR6A7erK9TDInlm6zg5iqgOPzu2ee+a7M3uVY2P2UG2Nov3
O2Nl/iFmCBFPJpRRZn1GgHwbgWUi57cBE8rK8ETmV7DrhuKKGSw6DYaC3VTLrhb/Zcybp+V6gteX
FUuI/wBQyAl/rKFP0+Mrixgzd3JOPEQyE4/RLZX6D08uH0JunUlUTx3O1JMC4pO0TDhn2TahCNjW
FBv/GeOcu4fe9Yi3bCoGtJe27rsL3FFaCM85nsz/B9tw4S9GdnCu4jE9Jg202d/gxwITkHQgHZLh
qtc6+ovn3I/fEm7pwmFRZ2DrgSJZTK6XBA/UhZGI+/sazRMF31LiR6avDoV2MCklSSMJpdo68OT5
YLQ+yFH614HSDFGn/FK/x8g78nAFlRP8QZCZABPOX11JWoE+fmJn9wgPsmOklhohwRq20WGOyUiN
DeWcntalrZ8NI8pmd3T3sEIb0dGmWFzu3Wx0uo1TaDjDs8JG71cM48JXdkBrbULhI2C84ECV1OVu
02CJdIbS/VZ7VE2MBnxb1mjw17Iz+KgaA6Iyd6axHYUKCMqyMa0rrbqsFiHS7Gl1AfS6W7uwd90P
KymeyHgz9MOJ5MkHQj/1v9yAP8Qz4r9UhOciS7g/AKT3XOeKHst9PsYg9S/4CSBlvp92Np8MfEaA
ECMPEw4qaK7CAwuWicBDhEaoYMG8x/PGORIFXHObl61I7Mnkyc+GWrfnxNh8CZ6BWjFt18GpKz3M
sVOHjgalpBA3mJeaCG9c+Lkj6fpy/4+4GzR3kqZmvpYNkSQCkHczMbHG73ciNhpoPVmGYxebBuQd
7PfV0AkuX+BU1aBpL8Z9/WkAZ4BUaLwmGN0ur+9asOFebtXTyAaKLBwJxFfZ/Fq/QvUAMeWcZ237
twwibyoyob3BB7TMr6onVGHyHqoZRRWr9hmYHGQ4euLT/4KkhoCX55591bO3HmJ3GyRl3/SW1l9Q
TDeAUh67hXIoo4JRauZdlkT8ucGaTSFtl/L+9uSgJZlqJ64jydEO6568rtQMlL1/+PWdCYaO1iO8
YGPgkkiy5Db2a5C2u/lLg3bMEUpzrJgYKvFP51/gGyPyrrDLeAq4KDe4pCGFEf+6ujwYwT5pvXwc
vkpG7B8rmO2N53sudmqXpSUngaaGFuJJ5Ozgt9lgjBrHvuxN6nSO+jCv5U61ObDa8yiZpKIgp638
MjQF0C6kZOBNI38CXAuWqe9mmM3+Hywgvpjug6zPYpBLhUoHyKD6e36B5RVqR3A2MzEhRnJh6S0U
If34SMpD8DszWW7sVVvaPcoSGC96I1cXydgtiabw5MQt3TcIqNEL3JNFJXFX1lkBftb6Wf3zj8Lj
YAuGAj8EsTsAHAjLVWy/cA9S5UjhV4/2ZNkhxdPmZeBoMtMxjWfvaTo/pJLivqPPEiYNdaHfoflD
57hXT7hAR2I8hEiCB1jWwzZPFX4c34C2OhwUnJMGH9aPctssPaQzlzTgr4ML0hvpSH/mgq9W7Qsu
8iwEkiSSGAv2iUlCzY/D7auLdon2v7j5cCQWMmWKPPVrRIt/Zsa03UxXPrxWaNANJxVHfW1TIqnE
9lqG3DKHwNV1XLLHOFNmWsX8VXfjSxu4ZFGgv0L7nt5b0gXGyruCeOScx2MoNcP/GBgMuB22zspU
4nTxrdNayq2LuK8cbE81XkYqNgnzBxNQl0b7VNMfvInf7jsEq93VYLJktTdqCxYwiul6vrTbwsO8
wUfuwgVNRhWCVl5LwTgLmC9Kxlpp5B9MHHwPBrhq1xe6+7MB+mnKgFRkQykx5Ozh61zYiyOLnSTl
3C6cH8RYQIM+TdiSbDMdikppDZTQWXvE5xxjkLFv8CS8zxTM8oaudH2JOVsct69bY/+DdATqg5Xk
Y0WnJTfY7xKHpdu4TadhMzX93/Z60vG7hgM7D6Fj3SJnQhkckDxXOcirSygwQBLKSugIczIe1R3q
5/nS8UjaIQr4zhh9rNilMZJPt+SJS74zUCAA4fkBguyEDdePbfMe1UJ6AWs+urmZCk9+g4s/4TyC
IIGv5vCellSWYDs5t3pRzTIRavXqNWz+4kI8g88STn1mWSGpuHKjxB/aGlCQzYtZofr/r0klcg85
X6kz7P0Ong5rxGwexwEgU1kw823Vey+7GPOBbqNGdPwts+kHr19bkzEajw6UCpN4WzrcsFZpwQzy
ijqhusWxbNcZTj92H/mMumjVNQId4UPFG9m7tL3nYiB7IYSbGrRZOJwSbW3RzedQu8KSzwWPhOdw
U60oBelrrC4Z50bZMIrrVVjHu/3t6K69p+14fMrK2s0ea/p13seugzjpuAeS2ZPuVuf96GAxzNrn
lSnaJQgIfQVcaE9jOlFk7odIMLN987qlLLrzsUbko9LjFQDTUQsAtLH74HEuNgdvT+2qSQ8hEdY4
rE9878jcHaGeQR2D1PS9RDZwVKa/pVNUDmsSVkADptDrC+T75QNuQXXAMcrpADMzJZO/cCP1z1x/
s32ymevJzU38G/2jlRUl/VsN94M5wvzg81JMeDhlbF3tX9T/uREDkACO6L6zUK77hM61kWw5nOo4
ECl2xBa6Nwpl/Xu9PljqdlQWO/N/HnYuvNCn8mtook69nwzeGRBkJLCA2ZyKYNT5KeQzIta7sGU9
1+dXqpfnhTm2qaxzfYkWun4pwm8Gs1iBp7gpbfcj+yrTmOgrlxKc3goQUSoz698s47Y3tfTGnhE8
JEvGP2hsR+z37mBXc+qymu/XiDXkN9EC2sebasw8n4OeHEe8QB5g7+ns8J+HoTrRlokgLHJaWgVC
fTdemy4uegsA/96mQPLlNqdCy2Tfb6Gq50ka4kAQ6LLzPTscAYwb7xjEiy/buS4XeTg2x/BXi6DR
IBoEGhhzm1wfMxVcoFTsVAPSrKqzG5Ve3wNxmdsBsFVFQm2+bE7+KM8UrrKnFNxG8YZlpPna8u7F
ctt220OdNC5EYGlMRS5dAECeHb6h7cB9KxvJJWBT/rztAPFrrPE0fkf4ikX/l+JGoMWSdPbtsWGw
UB24RV/ZDT5iAglKQ8M+Eq6NGwFc/QBF1RKAdFkmRBpfH8OgCvvtI0gOqLos17CoAeHJQf5RMpgP
qvw4H/zGDS8k9iKE4WYklDtrFzVFuKzTIE1GdtJyrhcfqLtNXeoueNX8Xkm4oA9oWuol6HfuxrdE
nikq1zxrfse3JQwffQHWKymvdDlEj8e2AxSbkJ6wGVsAJJ+xPAxzBDCZRmTezm3xCHGNvUS6muCw
v1UJQnqhP9GKlk8tO3TNkeDNtfHoLTCAWCvw70ep3qluh37oZDW4909lfkoAwTUDrxaJr0jnIenJ
PS2O0gFQTTfgn+oQXVC4mxBGToN/KvvahdKkAfHDg32otLEYJxEy2BUVlXLd/7+SAOB2Qw2OW43n
E2OMGmUOi/gX8QCIbxcOkad5K4U4pswI4oQdSmYsYtg2D5X60nUVMaV32Olc2160k1c9izItdvGG
sDrRLw92iKjvBJVuS4kAosZWrfk2eK51NWTyd1kjOsDp+BZI1qQuafAp9rCsrkJN2/kmYq3MYJkt
5hw2EUsC/CDgvb3SCPNmq8j4NR1MxxaIJxbRCSCW6JYUFdN1RRCcfC+dYhw8Cj0bbA5sZTP8tD6Z
qyudTNVKDeL1yhdC1r9IChCCcHNqEKfobHGfch3WAipbe8XYubM6CqqS8uylDXT2RqSI5Iie2GbS
a9wkuBd6HMviX4t6xnRVqiSrCNgrM+t4M6+xbJLHgGb/2Ybg/9SGhvVowbZS3MW9QCRFNb504NgP
bnyaHL2Wo3o0cL7mNpbm5h2Y9J9Qh5tghwy6kurjtuaEw62VjGbDNAv10bCUdYrnKXJgQHyyMIeU
tJUVUKFk6byHvGz92Zz6QAK0XeOMbIioxXPPGYwEQy+xFNimRNsxNNMAIK9UoyJSc9xtIApIQ2s9
z3XobisJASAi9EU2iICSEnvlrMly7KW1TexeQKL/LaGlXjJ+2L8le9AnwdltyD66yZc+aeisejiH
AHPjD6gSkslGxkwhz0Urr7nSMJYQvLH5Vcj8nDOP89EMjsoEn1PxjfRND+CTTPiip/PXhq3sABDh
DdugU7l7Qou1HsAY0UY2H3OtgQdv9r2mzDIoLg/TkP2XqhSXBD4slKq6LaZVg0ACdgd5uOGkSyKy
65NSIMLiyowx7eqTT7reXXoz/WTJT2Iolg8s6RcJvv0NXenCVgEAkgklp2iMonrm7f48kAnIgkaf
zUoPvudvvLAFTM1Psbtp/3s1GmZjOiU4S9UrMVtq292UKWI2q5GPBkWxmyUjjvR5vB8nENUvEe/8
97PkMoeD0SE4Ej9erQGyO4avx1GrrmeFeg6RjqV995NrYVHtoMr1thGATrM+ux+YVVwrwfANDEZO
803Eb6HaA31A6KVf09/6LkCEkecDCycBPbM5hE9RKLukxWW1LUMt5p4zu9q1PYnf9T15dVDUoopi
jsTGW0TCmUUmJ9dKz3xYnMmSat6l4hU2n3B3hVA29bb5xnJ9dtaA4OUZqhgOGfYIg8bDRzfQc+SD
M/UHJN3nveE7kBCairVE0iLjZTyW0KqNfZi0W00jA4LoriPBzLVmVG2p2HnX3rvSZwHBxUOHl4tQ
58kFFUDL9ShoItMlhFodj2duqUaxS2t6iZqBVyrhMHsnipolv3dbkjCWxd8iuQEYTuzlwGenaJwx
fBuf/dAus+XqOmkFq9RuohqC069BMIparzWdXyrsEqJLuHCbPJl4X8aWgEK1wHPUEPSECZG1y6qF
0CQbmgXyHb8XkAkz8B64pHbR6R8g1ZuZmmfaqoZSIihjM0Act2C8Dn7x0DP/2yoO0UNubnVs1KfQ
uo6jj4TOjtdjjDKVAyHgJqnVa2z6x0R4fjUUv6JkOVMtqpyjYh7xv3LXcdJZLOxbZWFrLPI/TDpu
jr+w0dXjnEvFcxqV/zmj8W5uqBgeTv+fmrZQ3J0D/xwNHEU6sBgkiNYyDEgwhzcMQ4Ip+eZA/ZlI
MSUZ7F0QMkF/gqh7d3m9GvXuhVDPhvwxu7R5Bm1pg8JG6E5027QYwKVSJ3XzLwEyJHQZOtwU7knB
iJJdiBKhTibMs8ASDCUsTvAfjdu0FlJEMXf9+ZzQJdhEWw18whdULCQb0FkMUWG9DDzMiO0y7JxP
WSFeopb9nAMlCTuXRXducbtXd4r5laAYklztav1gB2t+gW9/ciPUaoCWfl2Bxo8ebJB7JyETonBj
YeWl1EMW3ZdL3n3EW+o6Fx/sRPkPMCYIbWiluIbBGFD8fNhfI5LOGDIB/s891WRn2q4g3XnjBN6n
kk/H1FqiFMfV8Df1miD9WhII5bYyAUheYfJDzY95lz8jI7Xwne59yFROoZGd8xV4ikdyvx+qvaPX
ys5kaYrs5vfW8tNZ+ctciZOcDsA/0jGf3jn+ex27XUMeD9dBDoOpelCFCsP1IF/tbHMb3SPnnTFP
rEKG/0W573DXuzSnBS+cg3Y1bNFRwCr/uGOdY9/j42JV9ixolRncY4KZuE974JthkjDRNgXD2tld
PW41A1zNAr3USJ1QgmbDnL7z8G/hjcQwAcz0pybOZ0JIXfu3lZQgsiN7JXzy1kFQ+vv8Y4NtdTzj
6RIYa+60kvIGN5viIdLy6QreIISCrGsHj95kc/ca8FoRpFczi05D1dSfC7hc71t4SxbwwaHM8+XL
5kMwNh7GzEU8vv9E/dy1fgbdazFfb6G6Fdv650i6NcQkU9y5UjG/czGou1hviygmex6PtaiSPvcd
LsVL5Qzwp8DL7+zOmUoMnY7p0DvOX1V+TXhiLSrmtGjbWdkf6kfnZTOTPnFVqSWwV41/kOBN5n+A
mwKe6lr3T73qaCSgnj/akvxm4IzOrwEfOjLDrSprRycTI7Whifx+wKXekZHXrSuz3WPmOXufsF5Z
hbjXSeNDobF+OcAlRxPeXPdrvu1OwtpzUcOENOqOmV2Z4Tlhwpx+2NX3vnC6BlLzQsLIGZeDucFp
eK/RqiuiymVFiTSKLnyLrEWovjGWjK3fqw+GwG3ETMuY0vkXpHbpM0oB5yB4NLsVxOsPNS/9QCgV
G9KZmf0VehfodVppS74b9sBXQwOEoefvUV76DXf4zFh9Kqzr71ppb03KT5zMdcpAsfB2lz1jd2i1
JB5hg/zcerHNo/aG5VTug1ApOOVuLHHaE6yRG/lC1UO0P5YfECp+fWG4xCDqg3SW9FZwM8x+BYPv
BQQdwVtG3KOJDDFRXy4y6CJULOI/9u8KqmabvxdK9BzaJIBYcAa55InGioxjkCXGYNg2z+0DW9hV
3DfC60zOFxryehaMUBrkZueD/dtGxZLa1Fxdl3gscTW76R50F778ZOVz6vkk5ggDbXGl+c22vHbr
5NekdVMa32HJi6kU+h7CYd7Gkt7+rjkny/17qEfon8w46SSniMDuvWfFWL+43RQBEvXTAmKU71W4
+K7N68Pk9ePQnjb15FaDlyuWRaykidLtSFLOom9wMfOdlHSuyai7r7tdQm8J1zp9mchFFoXW5ha/
PiU5KzwH66fJeK3oADZZuVujY9FRdh41UILa+RIPMh0q0dbdC9mnGlhDhn5U0hsxIJ9FANKyvjiw
uKirtAA/MPPHZW6Ctw+oX1oXerDOZSzhIncz574pHesClwPukfKo/3jcp4Z0zorRnaQQmBxRQttp
ck2Y/jxaDakARvD/2mLvuc++9kZGZ1a5WztAK/c08FsxTZj4ScFj0kKRSdEimmiontr10YEt4srh
6a15E7Usaj2hy5XAtGCINXISMNvpQjkLgqvX16h0IU1Hmh3Cjp7T8bvO7QQfYncrHaw5YNnFI7VB
zJgOyk7F3i6fpLddn4QOucCSato0pApb62LHavlg7nsV0ySo4ocHfv+Vck3/SavUCTI7fbIgwGgh
QlzMvgkoX2ggSiCXOEuV3sooC6GMf22kJzZS6aSRkKfhnKO1UVDmJUQ21d9XDhH1XpC9Oc1w8auW
kkhe5xqfG1Nq0B8oULOx5WecMH5sSvIW/K3Yul1ce4Z1WzCiHYuWqJYUMTQRsvZZCQSwbSBJpRGX
mfJ2wvCMolIbHQ6uwQUOUKeKzEVOrZwXJd4GQW391LRoRiqZryxzlT0cTdJne1EK1qPBQBAh5Tdg
hZRFGLIh0b5VQJ1DB/u2G5UIHFih7usguXag9e7virzB+tHz3qegAQDU2ysreuw441czxjtEYQDI
rwoC/9rZDNN/1i1+1br0FyD82CaMTyOda0nXkezZAthYYAZ4nDnayosvU4Bo4mM2fOdkb9gCeS5G
cdx4kXVqkYpbmJtn57IqjTSaqiIzGHwk/fdYOyOUR0lRnp5aJ8YwoEXFHubahLmL486rwDHzrWJM
EZX7HmqtJDMiEDqI9nb8ASLz+52LrVWwUBLKChumcpaQPfLPrjI+Ns+DiVK48VlEUNwiiBG7XZZl
fk6e+4jyr2fm36m/oLGwVFDYVRPPcr3hs4TEkQOMia8xwUnn8PaTaNd9Qe/uZaCUYfU90tl/sAXj
3rVCNqzpCtM+csI6KPq2cTSrmsfxob2nCReJEfzc/agH5k9/Z22enx3AFnb8247HQycfRWT4IrTD
ZKcGp7eMxh68Mbtb6wnUrv4Sy+kGGH3YLWQoq4GmoToXhBjg/fkmB7az9B4z6bMclM2bYZshcpH/
sI1AUEMZPnNik2Q+kA77vmjEZ4ndCzeWEzlyU7agIL4KsSXK+iclBGgjNu7i5hh0cR9bYg3Yt30f
YI5C6hgvthmbIFhb79prw5FpWNVJQm7TNS0/f7LeIhtb6z2Wgp0mIW0aJBiFOLOFNLxplh68ZWxY
TK/klRZ9IbN+72DrzBh7szsI61IOsPC6IKLC0DEB0f4huxY64NMRjj0J9EQ/jzKft7J9VfEffJyR
VYhIx+2+4aYXS9RIIYmdpLbcc2hAu97ZN9wmJvTvS7qMHMs2Pw0zsmLioNOV9iKJ9tZY3H1+iy3E
AMnmmajhtUUy7Miit0SxgP0WY1gWY9+2tL6F40opPO0FN2Bm+A9Gfpvy80tCdODH/Pefne3EWH52
10156QvLhS4Nxq6QekKNwb6qWQDPPTqfOI2nappWp7js0eBlVtSl/A27P/FMSyzt0ABsQ1EIeu2D
75bfXnJOqkLc/E5O2wmyrcSS9P2U4AGeuaAfEwGoFxsIZYHM1ctqjDMcl0tP+PtmguZPBV/r1kxq
QEEqfoHg1/e1F7z13S5uAQhvb8ZmUA3+ZL9kbzpz5T8PvM67L6tBxwVVtTvddSnf4SuM36uznitI
+Y0WTIsG578ZFWhLznOR9ip8RsTdXth1hSdzNQuauFzpVmzCZ3AhIo+W4ayWf8YbnzcXlzf4+ugF
KO4ddDcz8CJFZsh9v4cRPNaC1qgJ0hBgOGh3r/HlFpqr/CVuKRaZIX+PRGhKp0z3+n/rsX3Ixyvk
4Kzm+weeftl7uuN4MWOPHcZO2FXJ1ELXghPB/Egwzp1oI9ah4lNHNrTUwGlYr6oaWtw0FlV0l5P4
aHUL/gaqh6mXk2yoj2MLSTiLTPWeXg8xBADZInX7OhJk5LHiQBtLLsfaV59JIX/2rfn3kpEEVQ1W
y8qAnVSgxpjCc7j7/+3iowPi4APNTONR3HdKOFjYIM5EtT5/hoWssNJSqO4rSH/iRxVJ7WIpReL9
Ecr4U65XTEv/dTgKvkzYrBkSQHJ+DKCfgmreII2vGeapRqOK6kSjf8WOVckG5uPr1ZoOV3q7LPKn
+M1y5KHD1LFTc74nbZKAioLE8LsNBKBMTRLwYvSpyEWSZ9NrTGeYFo1OLq1pwautWvK2x5U8wkzL
qUXV0nrHfwdhEbPYlTcf8213p2w/FbbkDWTJQKsgFwsbuR/Ir24W1sIkooLHTpIkmkf1ZDuo3uYo
x/+mnVTVrTOGErdcBf3EksqTEJ+/y14qDnWqGyrT9lGEt7XFVOYCpQQoagg40wwa1BVnwcc7AELp
qnkgGx688bOpgcBVmSJBGkX0EUY0kFlC/Q6K+NZA5Au032MXdKf2X+ehQnG82LOSxlUVWbhdGl5Q
8R7Ds53oyVj81izVQEolne5iWnbCIJZGajInZc1RfzZqS4WcbCHVRjptXls9yWCa13l5YKb5koCc
oMQaB/Z2VxKK85Lg69NPz0eVne99bwZsTTEJqXy0yII0KZoEw0IeLOxSc/46yJImrFNaQMdAMfUW
32E8s28QD49cFJh4sBwQIbP3BkSTIZ9ttpMVS0HtnCOA5yCqQ0DNI2mJMUG7JXionCQkzE2jn+1H
a+oJ7ewsdLO5iDkBa51tOHHuwb1N5dgd3kavAFwxZbfhVutQ5bPkpqEe5uEUvKoBMH1xxxeMp8JL
kzJaqzGIPsZGf5TTS4nvDSuu2gN2mh9PUIeYD6noDSYI6oR+5oDyTSyziZmNYJuKX7+8mgNXkO4f
XQdP65bGBEJlY0Yz8k7irQy8L5G0etWnRmTMBTMZKvy0vaBBQeWe4c22X/aEaf7Jes0TSUlgHxIs
MchEQAc9+V2hd1/XI8vejfbeYQy3yGnve8PkcEvJch3D+hxhi4LnWamOkneN3GtojiFSKVcPJKdz
4681xdgJC/8nJYi6m06dan26gBBCNNBqXUK/b1ypzreqCwhD0bkWqyNTpqMZ8vEvLjhDw07V8T89
hid582FgfCpE2D+mN+XtYTF81jD4ljJAhARn47MuOMXPOhT5pSeETsqOTpGFCFL4g1ipieUo8fqg
ljOVxr2tJeQbHtCuMbvaHXdgAmvm5/WtesZG623+i0CHmGmSlwOijM0wZmrOU+DqoQEP64S9Dg7Q
rJ+ov/yvA/PJoK1wN7FkfZ3DIo5TkC72ZOf6/4TlzSkkMSOe3kL9kPx9n1g3oAFcZ2yjAu3XKGtf
oeE/bJwHZkIcb6uGD/BS/Z8seFlNZKxwul7H8NMx1Eez3TcsXy73sLvGHiwBDYRDHrZjCaqLuZiO
bsTgOwR7OPey4c9l+f/h0b/4Chh5mVQxa5biDhvSjCLmAhRiU+0g/8/uI5PKkwpDq87glK7NQ7tL
nsGk8k9R3N695c5Xg9wxsyP+kITITMjiX0WjRgARJBZao/6utsGI4BcczJjAql54uuSiDNX0gtg/
jdR23MvU7T26J9qPLdFlxZE9XIve0SBomP4JvC+aC2NhLbzg9aoj5S5nqVWcw+ah0zwzYrG7e/52
uZNi8lq898QeTmoTJDgQBAstgxO77GHW0QD4jmY57MKdHwjDYyi4wWZirhwpDdpcPURjQHhziUAx
NIquxI58y5hgXEGGKKk3FHcraUGbgr2xb3ibFkhFl0Q0+wqS9RsMJM07L9ijEcFQwgmZGgMFvcSQ
W61P8wlqLwxiC5CFVF1ylIklcMpURQOK6a9l1Re0GZFW+VDhwgqQLmuBJ9BwQQljMibZG75vFkGP
uKm/rJCiTfOurTnUeJXZmuu6ZnVsXuVzT+OkrfWpw9Y8Y6tSdPn8z0cWb5Nic1BUR4nSxrCl7K/s
xtIXsu8prEf286srL7fY58LDNU0xLjpW8JZuMhm93X6a1PLgW0eobtwUa2cyQbcfc6jZXi17wjeO
2n3dt5koR7OJynQ2z9VtlxNhVKeam3wRzIV0e4AGQX+gpH4vxXbwjb6rALLH4SWX7jpctsfR0lhe
G7N9fIZdQ+sxcBNlEO6kBOrlPqJRiAOdPhWn9cRrKIE8HFKgEB0uVTRPREjkkiJFdtl1/7HadBYF
IN2VvK93EQ7Puf8j45FmhiOwbapRnAh1ZlUmiGllpuFKTSV6BPTwXvrB9vxmFJBkUyKeV7eeAj4e
B7udDVll4ROqYPep4pSJmPu+a5DyK4Wur/X33asc6qze2pHWB0+4kWarYROjp1FIPy/oSrUDd6Du
oLERPsFe+ZBEPIukV0UsXqUqjv6hxLnE2E2x1q+zsDfaJIX3BasEL9HOtLbulOmCDbETE+fTBThN
pIDajvlRyHgY3PA0okgkxRkDQDLFDZnhIEtdRtwjhLkqsz+0xRaV4vwXkmTCeoP2YdtihupDcxG7
4EtQysmgNDsx0Qsiko9nDqSdkIpZwktqlpwNSP7s60zsdefEZ58tV/ujxiRVHZUfL9WUyTO1f+LG
gNqjojuSlPfWkYKZGiN9ZrsfT7jAX98VDQ05DwrN+Bvw9GWHBS1y6hU7HAAI+YYx3/XmwziyMTnA
tHu3fRbc8G6Et5LVixZSfgcoqY7A5/hFluWmbHgtOkGs+iYbsJ2vIJc4ScjWmqyw8RYD5oOTOVEe
f6mJNFhFzFUdCPz90+NOheDieXSzGy6adHlR+brjSiviw4MDvVj630gyT1TqJfZPGFIbuZsWaMDz
sQYdpHcba6sdl3WKOC2VfxFA5BG+11KJGwWnNI6GNf3tjvrkJmsTkCvSiXQsvwhD3GXiQSb6qJac
zQ7NtEuG6sIbBlji1qycwHgFqe5qobw0Ctwm5UtbzY8fepDlnQwdJSwI5brAKJmMubbtc6PxTFZf
QSbF+k5SG7T1qyyjainXLfEya4IvGftPTX0i9GShL475UHOM9OQ37Jw8pGeG9RkGILyxlFjbPj/j
1NgqTgUm0CQSnTq0mAp2qLeGalHuuZaM45lt4qWfWc+W1k/W0ulWt4/U12mKeprvI8hGr6UKjIsy
j9GhULtS1IlaG6DZp1TlY7rbokiCP9sgIKvBnhRxpZ3qRNITQE3kLYCj0IYYwIdoYLzMBIo6konY
cAoxpRztoSYdM4YJ/f09oAUzHisAjcbs4dXk5nvCZ76tsAIeRYaspNSNpHh44w1KjkyBVvXEYdmJ
m23BhCTf6RM+abLvVbQDLjsrL2f/NBkp5NeUvoTEPhKP2LjftcYhwWvRVU+UzbUDOBfU8DLlny8N
tem/xKEIl+jAYkJr7sMI5ku9aVpHP0wdpqHB2n5ECYp4FA8+glWkU95wRseb9ZFUsHJPBbyPA95F
hao9tyFyClmxJ/3jwa5ZwzyN2iJLb+BqM/Z0U1jRJ5Buu7Hv/sOBJglhlDD2McEdMhAb0kIj8QLY
/HOFCyUGBylm/kAS0z9xNQ7eqJpatJSMUjUIDwhPtGmvZ+ol2NcYIPevsMLR5tKwPWa7EtBUxtio
P4yyRAmYgfgUfE4VRxPmmkzSJ06LkNXMCJ812iFsHzkYsJDSWe5W7N4m5hXpZeUym9/+IyVHhE1n
R4LXxsI3Yx7weYvGY92vXUT0ZuwxQhYCLb9rCmX6hifYiiHu0IK1ShrwuIV+Nba1b5tEH67uR7mw
/voITV9l8/HJ5l5XRns3b3/GhFaqJPTPc73JsJUVjF9nU5bXJekYHmEe/AJSr6brvHtKPrcEqFY8
BQOHLE5u7EUKA1wxrm7bQeAnib105bHc6RUz/xFRgHXHDEfmWjar1hZdr1KqkikAjetq63jf2CC3
ABeAFObX/i79nYrWtRUk34ZcCvs13YMWbMUTKC2Ml/KvhLQ4eflsQkkH90BvQZmyuYwupu0tWOPY
ybH68yY/dHo8jBSjFnVauEd+TdXa3DJxq6GC4Mvelg3jSI+4dVxVQ6Rez+4sOJjlCDX3i0w5noqj
/Nbk1dn2El8uSjZI/eea0g0pONR643++b46ARJsIOtS7QruCQsBcr2Mc0KCj1wwqM7PjSvCWzeMy
b1BQv+8UTXktyUcheWhi7GCcWPyXe8Yzwa21gyWjlnW/7CyHqM2fpJwEYuMU9/Mg3GlOQzpYP0Bn
vhko0p3T/VxQ7SNAu+cnuaaeJrm+S64UUA9EV/EErGKyS4NzNQCqrX5cKl3500uGJir+tGJH21Gj
GhhlVUQtjC7Z6p8u/bMSCBIx/NjIlLgHlF0icS1UuQ4b8iCnf67JcXsw/kJZVasGojOELsZb0o7F
Rn6hLm4fRJbNMoQJPFpbFxhJW/tRwdfg63E5jftqQHo3qzXnX4L5hySHPGtPEy5YrbqHfwdd1NCm
0Vyeqj7Gik0+xosqH3X/0wLN8dDES6x1JxLv9pMC3r/HB77ZUZ/s4apRAs6nfvJmX6AF1RiDiQRa
a/MqTm3nHYgW4g/9PnQQCQBuvm/+MQ3U3zQX+uafijlzXjDbIDdfipg0tl0DF9/5QiToJUdCkrlE
GggiWPr6QTqIfyYzUJmNthR2S9kkyHb4FA0qULDT8Ul2W3SAIswNE+++pIt7TzdZ3tqlItP+f0nk
GGvk/5ffyNkuZfIUiNxCeLc1IbpEhIJZG4+1SnaiP8YnujBk1z5fTM1y7vm4NCLu1MTPqILet9Z1
9CptPj+tKsEvtSO8eXD9ftOPFuzztF0jVN49zVM4utbcUJdXj8+nxAC4QQwMBbfx1ePW1CKvbMzA
yJkqRdzezmPEJwgncM/RKFXzkpAxDHbL++3demGweT0y3UEp2A26prNs2NNb5pP9JSfwD7/zRzud
Yk8g56KSdlzHqxofkWea3p8lTNLMavU7E8Ue9FcPCRP+kUo56mAQrJGKL082G+TKr5e4TcGxyVub
WIiYisw1CQa6dMyLQHOK9E9pNILgsG000/F5bBCh7bXUir5+3LQLiLwBwcY+f7+OOjEdUygDIiA6
wWpkB+cJo0wIB2K4Bi1czu/KvuTdREoadUj9RS3Wg3XrUtQ4o4iIaVmh6RxnoRoM3yY+Xy5KAHRD
lWZkx0mCbSABYbNci9nNrayoP06XF60FZZjQI5d1r+8qqBEH4lgTH4yDOxZyHfnafxucmSLlo6Af
oa4gV51c89/qgCGhLvlICrlqo3TRG97Dm6qQBvdcb/No51tyJ7ee2a5Zk2KWDJ9a1oim4GGhBJDF
AGCyf5lrb732HbNwP/Nz+iTup6EpjEkh21O03lkSI1hlPfbwGzhM3/ijWbhNFPahRcr3XpKBBAXr
n9ZVDl4v8I0pTlDqOyzxxow+LRB+kQWkUGKfa6MLsc8UAhj0SRj9uSziaXbAQMPYt1aaSaL6hdIb
/uKYXyOIhJsvi1WUbENC6GnCV1ONAWMpAoXMnMrvw60RyF0tgQ1r0wtWkbPzTSt/W8BN6abN/12z
Cs+IM2+y6VFQ2MxgBRlpLGMCfE2KJWjLJ/uSzUvNhGZLCwTGSAS42ybOZJEJmVYt56yvfPUCNfwB
/DyyzwasbVK/rfyslQLw2kUyq6ZSKKFykUCRFJAv7vsPSjFhWa0SUHN6/EbAgTiPndaDKMuB5/Q/
aMHVRiZsPbn00WRdI1wK4T5Rrz9iIulav1cdPBblfRGdcGYy4Y2qRcuhTWJXntBIoGnpz6WxCbI6
KAAgUr1dhFDYGeyUtX+mNTe3SEf8/rTNmXrQ9RYYkHFwzgwl5rVuMezFguVdXbsqNvv3QludwsqQ
/w6apJT11y6hm0SIZLH035/NoxDlekgsVLA2gA6BOyQ1HLaBdI0uTURXmXgtmLpCbD0DKuNDg9Kw
pzdCPSX9I5a78AV0+w1djt96YBrbmYjCxcqKNrfy+A8ggE64cuF4KiLhJXbXGqdGq8zT92SyA4WM
mC1FYvi0+ATh5Q1x+P5cP12Jwrtq26OeD+XSkeKp/gSQyFyj1hKR/Rq+NdBA8sj+5c6TxFbmmibp
aLoDTmkXD+7EregTtDzi8qLFR+HjXZVIHcXrUysLpnTB3ENpSuI2o2mnAIIa/bgRiRHz2scWeyY2
VOkE43dGak2EdP9TL9FlHbsMY9v6n8VZlcPzbPqtd9r8l62u5qzoXkyxf26lleynvTZJN18Tssh/
zzLdwXesUHGplNzBGcSD5T8LmMXlCm4lZA9o0L3a8Z7CgcQvT1pjbnr5IQ4aOCUi7MS2aUQTPpQS
5q/9Yi33fGEmzj4MexvpTUmRBRzT9Cf7BiXE8PBPBSpRk43kAxc29K57qS36xK9YbfJHjj2IVSbZ
6cM/QnWJzH9i0RYQO+Rv494ppu2MofDuy+CoaPdFr4a1AFzDcVsvk3DlcQSCpalR58HGL4npVGBf
KzBu4aVnjO6AfJSlAl2l2FgX63lQ6KJAH/Eu8VXEVN293w2TNEHkqFDTYNXKXlhE3Sv8vVQdaWJb
KeV6SDWm+CzoY0hJurj4JyRyEpMZieWo5tmJ9ozJrY8hTFNeO7aZRhNfajlroXVxuluLf9bQ5Oks
i13GEfuHxPaEgBvChcHPhe1VCzRCk/rdSMMFU7CsiNu77R8UzFkA974mIpJk5pkQqOhyjGgdmQ7Y
833AJutVuamWrwdH+qv+blLHUYS3gMIBWuRdtJ9S8rAJYi2NmPTk7nI2iGVrLZsvl4rGMjAgwT8T
IZWvo2coRP5/Fjyk1NqcR0wB7pVZcuV2sVYG6DimNVNGyeIUGhlKO70tdqMH1pZgEajKUlA+tiOj
U8IS9E5DKi3tJRU/DMXXVj9oJvCMmZ/HMse+OhSiZTDxm7y9CRtBX+VpWxcZFgjN+//d2afoR9ul
3wH4ntw1xJuF/7bKdd6+HIOJ3mi4IIjRwRIqL1yuPXuqzIIuVTujRnoUwyTlC1PHrr81dTmKuYu9
68pUzJE2cAbm1+OFqo0SYFN2fpp+499Rp94D0YigzYWizNiwwEB7RtLfRbgS4fFnVsEP5OIP4rwa
meo5fKqQAUvTkdzsy9UTHkQ+IkqWeuRBMxf6iCo4wI0KFgcGzEg77/f9ebq5MjAjQYUlnt/6VZB1
/exh0x4f3PmgGTM8bSo5xpWO38zioYwCjqeWustB9u8x2EeV1Y07R0Sic4ZHPuD3KMMOv/JzV9q+
2Lj3qCi+LxgMk8RfC0eHV0Nzj9WmzoXRInTZ8VqTqAGEsRkofpkh3xHxTv9iEJKjG1lUibQ7IdQ8
Rio907ODavoDnZFCl6jY/+u6dpDuV/IBqJ37oXjfQdTzPYb1gFZdwnVlMoMaGjDgPZJq2bQPlm+H
rL7rKTe8OwzrwOVNa0Drfw9ofWBzxy0Rvh2o7a8Jwxkf7E1JzEysM6xL+Vp9I8ceO3fcg8q2xWfH
Ur7xqNY71l2x3uO4+9S8Bp1ZcoptRUssei6xwtGEIbGKREF+qLUhk5bXz8RP/ttaUE+NrSTGZmUx
Zjk+sBYLWtoQqGHN3y+boRdx5MYSZ9CczJvmRIhWH1TpOGUyXZKYS39ACE/vXXEhr13FFuZlgSbF
QSD7zDeDXMTHKYZv72xaQKKG2szjVr3FRpH6ouuIHgVO24kDVRR6xoEnfJVpEJ8/TQF8wK2HmKLk
ugcTQZDqRphijH26c21/6EtMFF+iwvdFxGz58n/Cbe/xPetdZ+rprSGx3NKreLX7mSU+scNJUaVa
QqanzpPGeEfJ0sv8WLU0cAQ+29NuWEgns6XmlQt3wnzJmLpguokJTsfkRQg2PNqF0tIoj8ooiLpK
idXc7m4usp07+C+QQGjxBEEv+OVnlC9q1mEqa3cu9ZKPNZC557NsVMBf1Ox9e9TB8eiPl0ZH+FPZ
4jbb431v0sRfrvE7wLrt1ISo4QoGxRWCKHyTQK8R8fXzOi3Svv/MW2pZbzgNcEMhQE4MfIIgPv0P
g9qzix9cXTX1yesK3eajADe3vp4+NmgWei9heKEiLXtBXkemmk6w1BWmJnb4k0oCrSnak0DG/XZS
5ai8bjm7rJDI+3RIMgwP6WDkaxJC2cP94Oi+myMm1DBzaaTzoKXknI7cSmc22APv+NKRswiqnyPg
gNltE08myN1HitEhu11jyDPxlvah6Me8/lHAFl785rjee17Yy0wrjhurgLa9Ledm7gSQxDrhgdoV
z1jEt9RRv3Wy/JFDdqIveShVfqhwW/4mbtFRlqNoblvJ+rJaMfuJY8ursEDAIFnEK9ws2ZFJLo9D
LzvkhElo4dr30zxrZ1WVVGXdtzrxutOUlnVorEmwUYiPe7UoCco3vum0izSc0b2sAwP+W9EsOYsz
DBKHC523tf2ti4AYlt1yGaGNRFXZuanLzaYsp6fAFuIjVvuh/5mJVNqHSHvrZ2EGo+adPib7ycAF
FGpyaawTapU5QhtSwjis44slgEc1Dgu1pp+SVEAr2EtR/A/ZvlfRx6dN+82tEFg0CWFpb8izGY8/
uUDw8WupsrFmn2iCtPuiNoyTLOeMNSvBTyabYiWJsCMfavjaQE1L4hjkVhV6BXPOtYTFWBAl5vZ/
FCQFoniSQ4ecXSwUr6jpTNtmw+JkPsnHDZi9VX0D+m9270vSip+6jo14KktpMKHAwcVgImlVnVA9
y4wwYRTdaUViX/M+8RVqgFa5dbe6OSix+sJBwnv5iW6I3h+ow5PK9H3N0ZaY79XZjavzTNs9E28h
JvCniZ4bEuS4WBpsJreMAW52a79F1hM5tsFfPySFOXaJZRMRueU01F5jcjED+JZzbvl4mOL2ICIv
0N/y4iuDRRs+hOzpZcyiqiHDdUrH4U4z2t5+xnhUEQgE2R1Q1zlE4QvvfXogtY9UWb4zHzeT9mFV
s39A1jp/B3UMLIeJZC13+wMy6pe2v8nPhQlPuHfAzRHqUqa4+8m9nZSuIsCKZkWtQvQq6k8+iRim
VoSeqOEZw+TWTijoDtAMVnZecGsSWSJ+jKN9KTvUKEHW6H6JV1+S+mYKn/WvZVPHQsnOQ4Z4T0q1
EJ+Vkb+HkMtVhpQo2xOI8R5eD46xZy2ztKLUe3v41Iju/dx+MzRiOQgKt3XFyS7MA01jl0HiVse1
Mue1bhFLW5ATixUG9lWG9aRHsfNE9LMgzSsK/n5RDI5ENLHSDuf0lxdBt8lILzantKJjkYmAqq+j
YX+yyDC0V/HOOFEWdpMhikA4JeICN8tvUoaE/Vnr6AC/EGtNgw/JCDwJT4rdt+Xbe0c48D0pQzC1
OudMCtuY6WahgHK016G2zDYMWDpbOWlq0y84gW4jdbJtaAJv59ubWTOiFe9E/717L3PBFVd4NfZY
rUVj3pYwFK+kJqXdQVvjdYyNDTw0Y9VMJ1jKcHqZu6KZ+mXbwpegdmFof73+XXM/R3fmXhB105Nl
c2L1jkVt5Ad3nXtVIvTo3nHvNXBGBrzmAwKOxEoow7Smc3YSgB+GoY2Nnv+PAMHw/DAqkf8Dq5rv
QfcbUQgKBuD9rYmDaEcFk1EnKfzg3oVwvCQ9pOAQH6uST+SCZBZMxRR1VDadE6M4BBCOpJTx7TwU
lI+JzQbfFxe+kJHKLUFLdY7rBkWa8bFodTPgM1MmPb1LkxnXaA/kWmg8kf/jB2P6W4W5353s9fsC
rlLb9OOSKjUXjoNzJgUITmNxYL49XD+RBDD5rT/T0f6WSV+Lh9ihzdVFsh42MttGQznZ5eness1E
WNQ+V2xZ2cx3AeXLXTwco5VF/A64VYXuX5s5uNLYJ3XUe2YZsAgSYALvSzMdMVjAJa5fyS+ZfB4C
EeDb4CMsviYCWzN0dspMA7eTDX44rkT6ieL1XfpCgW9gder/oQ+fPpfM0Fk027L7rv0mYliUACdN
8GZAcf5evarmVKQ+ceVBoNRrkHgSDRyUlTROM0TmbtnU8VRK7u9uDs4mQkMl/k5RYOctpIIgWzLk
bIoYZRns2/bj4BiF7kh9sT+Lse32bEKe3kDF/o0vA2tFjgMBq/a3Ua/Eoq2BNnHLjQ+vBB4iOJMv
0H0jkvvC80OdDmlhXZWIecW4A66Jcunjb6knYbznxoon0FuHvh8znorLE6pCRNLiv3wzkDpEMF0N
mmUb7R3ai5g1obqDH3SRLlQs1ZLUBEA9xCMlIdIu9hB1RTJhflGKAUqQ6mx7sbD3ihZN+KQnZiMS
DguT0UR3QpAFte37fAkhvM8HtBQoG33fJfgEyS9vI1u7o2oG6qyPoiZG2lrGQYUpWXjhl7t5voQz
LzdGrjWDDNzr1Zl73cix6Vmz5dKN47P9BpHJ6w21ijYAHvuchaH/QE9hR5O9PgnLah29E78jKdty
6hI7RPR0Cftah3ncNdGpj4hmb97PM+oNXOZ0RiAahrYdRIsbJfs5HMiifpOUZfF1l4e1hdOavF1s
8gCBTakHFOxmzAth/wUHCX30fha/pbytRD37OEajPb3roK87dXMm6Hgv9j8tgDg2cBM8DE38WOmk
0052VtWfZn3ZWOd7M/WlDMPzj0ImzAE+lx3BAmXSldtY7by1LsyeNNveN6B/cbOe4DNavZFE2Sxv
fO07jP0ziBaFP+5pCyaFVJhQGWa/StmhsGQznXhmPetmMfoaMkFy298xwR3nfv2MfYsS1PyO8JBy
jAetBkybtVEE44oXpwupeOogB7MjXFxTR71hU/AlEWXH/FFlj7XTerQIXyZs0Sf6J9ha1arIVqtz
oMkBp5aiCqqnZS8vOM4HGpHx4E/nOohGdNGrU92GNtShLSPZQ0EgG62yFNGJIrhAQwNsA0NFqUeA
wgAdcJmtaqYPkD16MRFO0Qpt75YLv89ZYWzjE9yzlsv72oet5WYpaGhS9LdQpBOyQzjuEQkopXIs
kTN+zIo5bApbaLG791hPsmAgSZTG89TxNcAR3Z/J7lnIXkS4toI7OIF7/ecIoa2KLSIVxvTj5T2M
73gB1cuRS0MdkHppYh4KDJA5rsHg/sOwcVk3Adna6yMM9uLyUQ0kAu2wHIqNV1TzpBbY9Axk8fkY
z6/+zx26cRthG3pOTdst1mJaa8q+JkwdEIHIzfUtfvjY6q3O7kCpFj6pG2epqQOGa5kJvwRlcl7h
nFiDYYqFH0wY+b1v7+5E5pqK8CemdpEqd9oJcSpdO3sAcqueaHoZyM1cS9FpTlsmsBK8GzkG+iZp
3/OJIclMYD9XbfAPYyBIcQzld28YCZKeiZfjGpWE3LotoWvUDOuokJKB5Vavc0xCIqTBYxbECSYv
g3/LSkx4cEjJK3BfpiORzvNHrIX91ZeLam5Wyf1rkQ/0u4wTGHVF4CzeLwJbkS1AdQ0bvm5CoKXH
+3oh5EgJbglyqqWoo5rVZsE4WQJwqTEVjEE4wPt6d0KtaXf9CnhRCNUL+u6KN3170/C2oAwY9IGk
pNBO1cFG08XAuxJkX82fLzih/RDXQSEwGqeBlpEN0B+m62y4Pkyd/1Q/FNI8fLTH4uAIdm7sDETH
taj4+jk4WBd6NwmUGOvTjUNdPbi5K2lzGu4+SygdW4g6IOM86g9u2vbjAvY9MBq1adRugQqt9A89
JLlEgPFI/4uEcBr5QSPJK+HoLuIn9UTqAkdPj2roH0HI//jx7Qa1gAb6mgQtXjG2kq1P+jQLXso5
OUwHvsKijS8ENhNyVE8GC3I2TmI0yWuMlDE0eW7G/1N2PLsnqm9jX5Nm9nA2cZCKOniYkQSZvGuS
mzxWUFOFfj5D84x0eNhNk7XK/pFbmeeGlgs2YErNL2K4vh3yfx7+BdMqjWO+b+zVlu/14qTZ8JAS
9yZVTjUvd4QB3ubIK586aSKWmpEQSColXfLXQNXDpm8+JQKQcQMqG6F5LDtFdxIH65Bg9qJKr0H3
36BR6yGmoJK2GXMUkcrei8qjVYr/07zRo2zh9Wn3fLOCSdvGEbyu+p8or7HnI+bnnWzjkEXydl5l
6OwgcEqiwtqruKJq+ZemjylXunc5fmFC4J9IWhPefi/h3Rkh5ymQarhZzD+yXjjA3W04IvDhcdSa
Mlm8+CrZOEkYlPRlz/mCui+LFvOB8eduQW6EuI5NgK34QRV0UlhWqJt+fp8xrBTg2eb/K/EQLjQL
G1kY8gx2YEIRFIFuO7Zt/RxmPyoK6ME5MwatBmkDKLMsR+BZ9lVF29C4jtGmFb3YKJrHYvNN4ii0
sGvAHuM9lhetSl1z/SwGpi3jpYf8oPdBj5N9w3jrqUrp2s65lc+jBVCtQf6J1PBME88XuUE61BKi
+/YuZ2iyHbetgtQJjQPQEu992RCljVgsyZpSvj8wHhl/nGV3BK9tUcoO3+JIq8VJzfT4JTaapkR8
bkW9neCyyk6qn8l1owurQXPoTgvr/5antGlK349e0eBaoXpqf+2v/7yThS4UGme8sf83AbM9yuI0
S4bhrf4b/XScRMICoc6DmvhS3Z5q0HS8vV0UvizHIt/FQAYK/65107og09ExEgcCp7KQkN5ETgwx
VSRUDs+0fEAhdk2hRqJvzagLgFp/xPjd8QXzVtjmFUFVd+Y/adHq1y330BglAJ5iKHugeIi83ARd
lCOsSqkod02eEliQwJSxBFZDNBzwKvhna8bYY0E4fMl/4JrN3uTO7jmaFPPM/PTjUNhnwzwjQR+Z
7LiqbCXEZ0x+a1itwph+VgBEeLcUTQTwJBT1KdcMsDA6m+IMJhFSiHbt1uMDkpLpKu/3RmV3zFo2
vWtPPh3ctymGdU1asC5LaIKfrQTW6vDrBU3xu+AbpWsatpclOfypzIsC65bCSGXttzwjsd4I9p0T
nZYouOmuCIZmI0BST09lvSkkskT4MHF5W6vTxrUiW9sgjZSi772+gWDAED8yQhtWRlqx73FkxTu0
Sw0O+sdAJ/TA5rN2u6v03qBnJvrbIm2EzeVmRc3rLAAnBI5IPu2dD0wiaAt8tXEECj1NzSM7gSKk
ur0wK3Ijai3HfXE9EtWFUltWQGCcENZudGmqZce83vY01viwpWzurKMbatRmYjbyH9dSt51aFuqb
P0eeglIy5d9nWVWT7RAIPurvom/2Txfao/DIu7ZsXkqTRUs9WdahjEl9q0Ziuw2vqPWgehe4ceRI
aUF9RK3LYxSKvzZivd38xkO8cBIlQx/dpL8NFlKbYgUW4EhCNsh7DVVehzyvIU6hCw1U32d5V0Gf
nNwa1aUcqOeT1PCx+NhBCTW0AHUoG2ak8MmxmHF1mfFv6aJaw19SzaNNMNa+GE3kIb0hL8f1anO8
o+MomXtzyE1w8yAiwj3frAEvORTyo9mhv0s7ZoeeWmKaqfemY8cc4C7OxgMFw/68RZslY3o6U87Q
66scmyCm81aSueGGUz+8WmJi4cnxQcvmyfzJOktSHj4UUowc6TKxdAXePhSAReeDkOJStOEQe6lO
PGA/+5+xYDcfJm+lbhh4K/4hJK95mniKCTqomAPVioz5ZPZ7av5TA8ZTUx7EhauWZvtjqtkXatMf
ZjJBgHsX/7Oyu3dli5iuBTFdN/CMEwyhbFGZ4TzWzRZetvoCsBdnF+wOk37R6GDsKQUdpr3BFuwT
r8V5znT4AUKGEKEvX/eO4rZ56wfgWYyHBi1UAH23xmrRzukTQA0QY23fRT0h8EZEal8DtqUd0VlZ
MDYQbONvmJmvghDzeuvVGpj4RJeLWxF3qIHnTaSbEnoA7WHLhGqpSMsNbod9oRicC0YkuczOaiCg
QwuD22NfVTJsWloKXBmzTbiWW8+ydzxEUjlMQ80l991XCgATghq6a3Qo2GjHMbVKmjg0pThuBR4s
gl6eImbJ+DiI4OHrpFCJDmqf/ci4NQjEXknMrnR3sOkOCZi88YdAOw/HkBiMY5xnahzPO4llnEap
FdmE8xc1iSl7qAPUyPQ4atJwdXaHT2BjHH30bt+PMiJGTREIOE3KUg6qbZyuoGfBqQdLw2IYJwtb
SeLnb/Q6auBser8MzOTmOFF/BGFBaR+SVTln2IdhYoDw0tY94e72Z8hE9ompsdI0k915444GC8Oc
QPRenvmbGtqKYN4b2ZJMvK+fnueOJD5GO0S8XIK6PqS+0wDHiBWahSmS3Z6kYV9aYIUdNpv4ETfV
pWR5stVd7xGJVCgtxTubvuQbVXj4ot5IIyu0IDprrBIy2DMlR7shidSlKgf4VHYcRAVbI6bSY3M9
7nzgWinfndJ4tydWfLiNzX057xjE2THVwu7OMcrUTJimo0SINZ1//go/PFHG7rX8HBbiTd2JURnb
BS6YUSxOhieAc0QLqnqLWXZ7edJxEvzGt8SrQ43q1u5+gWRnUOag+CjBxZmQYMdCFefI1H+YPWUU
gK/mmKk9dcdQfQ03Kt+bH5zThKZi63oG+B9kcslzt/py1bELhZ95nxyUcwXFcXxAxjEBKXNNMcsr
fvS4jP/Kl3FhPpJYxID5144iZy69CPcFykTBWSLf+T8HgBShcVeG2xYq52xVkkj10WonFiSN7+k7
j1gxuViux7uNUFWDpHNZCfOpjEBphdFDETRQDFgE3deWolZ7eJCg144eYysL9X68K6zzBLqjwNGx
W1TXWOxxUihSj+L0aS/SoaH0SYJFkvkSWfLUVQ6JlczvbD/TipfBHm0g85ta15ndcU3q+XzeSczF
AauikdTgLvx//Pn14vtoX21FCJvIpU9lUyyMJKN2ATRS5Xmu0HnV2nVna3WYrzfMTDMdPhyW4I1I
sHqaGekX9xDvdxiLZTBvr/M+Km5naMcVJWEOVlzoAwAxNpJh/b8Rj7vtZi2qz7E9vQbv/ATQ/oqF
YO8NK+dhmlOUWW7WPxiIzz3RWIeHNVZoDjLwDODL/IUlugn9iFQjGeOSlpB48OZobwUTPIz4o2Bk
fX8Cn/GkeblV/HEMml8Lafd4AbfsXUy6L9yHsv7qotB9F7NnoHAhewHsxNkJtDm+RNCmmgs3XRrN
Ei+v1dpRbqoPGnXshw4h+kYrg9fnt+qme0zAX28MGxi1OwQJZezYW4O+JAnwuHraYoctSEm1bX2Y
kaJh1HJt25W5BarN/FtYqZi04yyPode8cy2ECgxb6Q8/QkQvGqXGVsOvzYNHLBtb8Yf+JMnvidop
N0g3w+lT/cY2YvKfRs5oW1VY70/HWg1XvqxpPucdFK0pnVk1QKE10rCGIEr9WNPRUqd/Nv6hXaVS
sAVnVsD3OWugvdZ6+mo18rXE6I66e6y35TWjliLPuN6pba+aN67dMFthwgdZ44KjTAtH+zCM8sMr
Pw89+m0mMZ0s/R9SovtXj7bzfsB0Af4Ll8h5FDzkUq9dJOl8+w54iRRCYBKo91bUHvAAUeeK/0WV
wWj+Tr4rAhnZOpeUbMn2eStgbkM5uWKw5ycW138W9QKk3muMYOQIdRJyE4/0Z5nRVeqSYDi7jIhW
gJqpmR5qiwMUJhknjacUb1nnt/YuRwDHqqx1UmqOsIF07l7C76O+hk4Kr/9bdibCi9BZbCHZopyE
/DrTkZ19PiDj/AzLzJWcVXZOBTLc3qvFG9S941I63WWY3G3HJPZ7cWFf2q0cIgdZLdBF+pkLE7sJ
zQvysGOCv21jOvP913xD10YAAnYjgTw3tohwxx7e0pX4/Qs5aHc+o8T8x3hVqXv8mMnLIaLWLaDV
QVpH8Dg8qBXcNFmX1lPnRuZ5wDd5QY+GF3DVT2zhOtfTaQ0RG+ZbqCr4fEfdLMrlsOHL72YyEoLd
HbpAN3ferql92zNLfSrOOURORfwcD/Wl7/goDftfr0Jd+T/USEyzSMqH/LieaLbFSkqlkr1Brq/z
j1sgW7g5FGPDfVf0QtaNKPTO+hSxVtJW9d7H1XmM9ps6+FWkAB2qxyornpO++1BMhFnclkH7km9w
LEyW8pNZnKaqMd82HrbUylsgAdlngFxQ4nx5ijVRvVFcrt4lgAR2rYPiqGcVgAqUAsWhveDev75V
RV5+odBdY4p1riYWRYklk3siYTyd79Kp95QoUxURJ4gqhEbgeRNJrBI7ya6PVYppi/Nc8Es377py
GzLQiuGNJJFKmY1tRKttN03F/8b/prgZ2Yon1DgUd8OR77wonUwZbgVYoCiqNB1LOe0JcX5ErMP4
4YSYoqTaML0Zj9CDzm0nv+4KD6igZAPUPWavLQG/lXLf/oG92h4nNVdC7puKkZhuhczciMR8cwkM
2pQGr7dR5HClxqRMQug/VNL5B62110F23uk67S6+atTqvCFKP+TgldHMHQDfmr4mw656hs2VEuif
ShkIWnkFYZKgAQjmtUBLlvOOsAeHy3Itp4PE3xFSu18d4zJ/bsMRtu8I8r9rpIPzmjFksqrGYri1
IUa5dOBcAdN1mgen65DCgbBVaVpUqX2zxnbzSeGygtl1k+MrxHlI6HU5orPbn66C8PUoAODYEfFq
pDpkLkcQcG16vwju1hjbCgwWdXcrjb0FnUBBWDiLgglAPHsmFNM7t8p3QCuXaYRdz5xgJ8Zb29cJ
a/sT3TCE96eevNuW0VPPDfxL7aqajq0qTvLxg+EsJq7q9BKBaA7Rk/hkcK95j9pY7NXuFnlAgaZO
zpiRQmCwfhHb+Ps16AhNaHJTZnODLuac/C7XbyVeEpKnGIl25m/RuqBhKpTcm/MGv60zZfiNuqR0
NgWFBtUcrXE21CY9IgPtIhnvxrFSpY89CwCXfj/g4dB7zhQsdMBoB4+scFTo0Hu5we6DamI7FHtI
Y8UMMOvXVpKYfGLwZnEFlg3u6zaNbNCKbYYvIww+vdNqZggqoTpyJWs5W2nKrvjVd5uvQbizTrBs
XLXSd7nR79khbKjsLBhLHZpgIyx9QXDm8mdL5jY32+4HGsu7ITxDLNYKP12KO+AXjguPFLZxE458
gEgiwxrFp4J8k3e3Xnj5RIP15oJPLjzmQcJIsQujtnTxn1wFJinfm/sO13oHZIzD9ABV6cBLbMV5
REBFsUqzadVyjMJd6yG8mWt1PwhaoeJNdgPlGXkQPSLra9GzdvjNyoqiV3HLkpEXQD2jllpceHSd
HciQXRNQXKnGn4bWWf23h5sd3+4DvsjjLf+bnNOyi58mhFxGBOvP0BCaS5g1i6ZTTt+bfmFBLXIz
lA83nMBcuczAjkL7DtuEZANOGnOQkXqyLY+ZWhs8hNMckiE26F4lWOg0qlfQfEozB8UcIQk1otL1
MyBqB8J2PL45kQna7mpz3E46N2IVD6xbG5Dd9vMv7ZDjWz0OfUnLUqJwY5JeUK/kSfkgUiPh/rkw
YEyljpBYPAkOTbVpvbWHFNtOf36VdPAGcq3L0mXDE2+VeTt3ms9X2OJncGZXrpt+ekxqslW0bquh
R6z5/P5ZPnDaXBU5j/mtn/uB7qXCMu2Cq7c/pbIs8/l+Z0KsovrIJH/swtgaC7WlERedS+5HT8fV
JuoI5nHqm7ChGQWH6E1Kf+jS72ci49e7rSxG2yOCKee+auofE7KNxB7UCV8ZufaZ5G77iauJSRLl
yi+0LcPOgsLdrK2ifelDGKQenJeNUu9yIAYlOQWoNt1TxGAVWaMZDDpWiexJCdZDdlWb+sFhGXAE
s/uOwoTXmyCDmAXDn9wi8Z7qOT/5AHWzP/kHTHO0Fw664f6tllSGuej6Kmi9bxGiTGKc8XinRxs0
aY4Jz5NA4gFmKzXGcg7eZwYXKk+v3Ynm8sWOBd6ZntAMhOBh2moh7+HZ5fgf/Lqm+mQjfTqL7ImJ
EEzu+t9tC79HmGAChuXjwtv6hZLvScFrQE+jrEeEPvnlHRGC/yiz0ZIpfzQA6NLCto51M3MxPLjp
KSunp7nvaW0wQIds9dx1OA+Qc4x+gJJrx/2dGDaIqwAO1Lug6F8Kj+F3LkcD2wChe69ItOZvGdaE
OXm0jm+xNXCZ3ooovIDqaoWNawRJB0lvYpRDenayJ0YgIIhboObvh+BB+/x9yUkvJ/Zxagb20tKS
2fQBjAoB2bkCIdbRENmMoF8x6fWuyKD5P2JtNi3SocUNEWy/yNeiX+/z5+m2QtnA69jdo808IqAE
vMeLGBI6hipGeI2wTPt6/Eg2SVf8P5h7K39SAukDufASEG7elQPWVGpPeyRDRqOOIJ1j1n2wmIxr
P+n4BOiPlsThJ/d8pmEzUc67d3poWOJt/GMkqjUXtbVRxkxwhSnXkeM0waGTsB4ofmyzkSGz1t46
PByaaW6E0pyK5nxugrs9pqlu3xOv54mItAu5OHjWPP/PFOdpnbWmYXYs5KLNhYMeUNZouoY1s28O
DCDUSpD2mWQDIQ88UR7JhSI/O8YVC6oNeSpzHOZr5hjG9X7GizpULINj2jn4DmPMn6d4AkV7cclH
NEry+Y1mcr5p5d/UzR+dMquCj9QVyfMPHbwbH/dQ0Mk295m6l1enLsWXcExlI/X/uFKy0Az+JQNR
VmfLikXiSWaofjw0ItODq5/Vu/WSYS/8+T6Qxls/RqevqN8wYlOJS9wEPibe0VGVwu1ubYxQbEGv
L3BCXXzGR8AdOTWD05UwnO9FLXwvV4WgWoB7ZAvWnTzhTGELGOK4iYXyZDDu9+U3CtZh2SD2HnTH
bykKB1vqFloo8AUcTnLwDUIEDO9fyu1kUUHIiwFupAaY0Tlfq5zmZ+glGtw80mISVQYZuPvEmxus
Z+s/x+TF/syfXBmDzvkVBcEOqZj7sLRwVUqdkCv1fZd84LcRnjYWpONGkO2PrWPeJjhESXAOJqP+
u3+5RCqNoGSCDGE8Ct7yzyE8JyS86OJvilErMyVTS8YEMZiEjX/iYs0Mm0KEl8oscj+8jSwzeYu8
e281QTuBKxzTfSGFokJzi7ErchnOVtJSqof6qsQV7yPktPtYM7ubsdnjRCcVbgC1r1UTTb7DMTkT
IPQlAA63J47830CmXA8bnIHLaoAP49v+xaReGzMHZ9b1KN748TRGYJ2/jPtxs+wAzIEWNCeJrF6I
B5MBaf/ahzN/embDDPCUXVikttGIDXuiOwS0BJVifSAzgUygzRmEXdQ+mSLnhof286JlDyRrikvj
b1JUe9xbCtSvSkVPk5WXCVGC9a4r6hwLOOTGjt8fdPUF/33f9zwW8DHiMXSq2jbeSdjUMNCHDX+p
YUDh6zcsNgxfJwK0Ng9pyvSYVndaLHjjjNJPLrjxyTRM9LXoqgO88IAZEIzBZNMXCby7/j+RIik3
PAUMmjGxmxkoSQG5A5BqKo6Jlzr4K5dHV2qVz2N9DSafmga1E8K6XfONMWm8tIoHQeFf6ZGMuYPb
NV15XSNdjXWgxOOH9qnD99GP8Rb9Yk/TqAmWj2f0H4OtKvkOSJJq9sqwqfVlFJAOQfqRfmnWZAek
rxntwzRV9F7JjuLal5zdcKYT+yAWFLlqzVAIgs0oRIVnn2dAZzNoHUIUdW4HZ7MtYr7m5OGThz3Q
f5BjHYnyij9N3hqfildEnOwVGQSULjAO6fskKW4nbzbdbav1ygtfm4EMv46ab85ZonMRkcQIDwGQ
i3SOnx/OsJJrsVFdk3G1+5igdDwh7OJICp6f1Bye128E0PqpEx3ffrpc26CZkfQeYKNeXITiqS3D
RYc7JwcRBVUWFMosg4EbSeA0MHBUSMnybUoHudvw4g/uN+V1aTpgzV9twLcO7RFh99tTxI5Kqy1K
brE1KobGHG+kVxCD+sP/DePGdvn99JezHBICgKTQNIHPluvgOsOQj9wa1TmwcXymV5Bxgi1tx9zD
esMcubHKNFmWm21WpMM6/68LXoR5XdqayLRvZ4pNXhkRoNS8QVfLbNdoqSAwnzC5ze7K0eX7lRQd
lYj2FZF7DtSkQnFYYgOqI2aRmxY6nMC6GZFnOXBOix+45pDHZ8Py1hy4YNY0Z8c4a6gGEA/nVzpA
nf+eBOHDiGiYCCbGIxnxjI/xE3BPwriARuTM+/qW/ao2tB2tUIXapWGJM3cY5rFBl8m9ayCVU84M
4pzM/XrpczD9t/o/kXcuGwn6+2uUdswJ0wa1o1HujXxfsx4D4pRuZu0YPcWS2D537ie4Gt8auqZr
4tYB4WZbeXb5GR6Z6rQqymgjZis+MoA0g6OXpDTx61eZb98C0SJSNcqVlYA0DoGut37nSmh/YaH9
8SU5BittIEeHIv2Q6yBRe9fGl+IMLQVqveJukedMqQAUnhWb6m8NgbjNvkqzOT92rbo/zydXbPQ2
TpbW1hMIs+geJJu3K/a/+WbczuSHNYbrCMJh25d1wg/j83YC744ZECyrvZqrw2b0ME8XgKvPoMB5
lWjETZZTYAjQXhKV/Wsw9BTJwEP+esJoWCCg+T5AjGhb3ngyDmwFX5fQRpu12G1ds/iMBCV46wye
rjMnS8yi1MsCYJGiO9zd6o+Kg382bKeKOTA7modEjBcYHZGSis/MTVDVuRvaDbgRdBFyvjza8xhk
zt67oyo/s+BfC8+PbTaozrmv+x+3GftrwdRiUux3mX1wrje1nB+w6sJBxby6mbosnm3v55Fp3vFs
I/ryTrDQsnDv+iDcEeXhPfpLzevPvRLZedpSODpeT/Fmd/F5ClvK/ugwlKo4fVgmjLssGb5gG89w
Yi4pFkKXC/4lVJcBaLvUIhuTrA+wjRzAWaE+0o/N4uMcyc0WMJYk8uw7AdzEBredDh45xDHdNHQ6
9cnoihUha3vYbbspCEyaHQjzHEP42+tGvy59jAIbyuetKrZW2vUvixaHxk9F6NnxycHDkwg7D9ur
3xeDXITKtlHG1N+LNW9Kan7Q3F+o3ooZj7oRlK9LZnQvM63fC8PQ5jihAE5/FbuhvhxyBRgklWsh
VG75ttDrovmYoU5SuOipdHCiWEO524vNiF7duf09u/IKYbYp95cImeAAdv/DvmLUkPYby1bC95dF
5/pAi9YB60prbJnQY+d8OyTU5l2Deu4sZmGPSoF2C3h+zhlVZ/h3izvAuZbiKySAZjZ3tnwGrJfV
QJXslVx7Gd4L9zmA/SI8B4/SCfATGTaTi6R4gfcpOHlRGc/QuvF5kqa38BufmdgLKcZR/5Klba5H
lHsg/edEVb8VYlIFb9YBAocvnV0BkbAbsbcK1WAuGFx877cHFiB3XOhSHfFMbzyMeQSPYNWAiALt
EZ4Te+Dd+jlVKRF0fcFYZeq5Bi9OhEt5+j718Pc4cEP8fL2uiyr2/E9noTWXfnhm3mG3rk/FGjax
tN8KnpfpkOk5T9H0ifhgk1nuu9XInODt/hvMSR6e08Yo3Ofag8Db67ptIFalm8Sb/lkaG4a14udr
7WjZ39lRFzTbwMMsmhfztr4Ogp/pTnzB17cyLrvgL1MWMCw46bh5z1N/IL9aKR0J/wcMzuPn0gdj
/Bd/9Cy6YSIRHRo0+3INDVfA97N9CjLWlgYigCwYZa+Wwn8nEg7Zet/FAKXdG2/SiTp0/TwkJBku
CLZtzhN+jrAzwkbfdiFzNKOMExElOUlWAjoxwZGM1D1knBAmXLXempioBjjbvq7IEYehUd89ib8o
/FLXv9brmxDukV0HPOhuRMgns3KUeRisZDfVuVMmybA90eaxi6fIdCBXRr4CjyNAfFB6b0EIgRbu
qjK/In7hBGxb6FWUvj7+RNpNX9hUQBLaM2G+Tv7uTuOpiO2ejEXfD90QuN2QPIAg/sef2n7NDIUp
Yd6RX1xsUEdW7lpvVgBqrTtaSdOP6ytuWPLLSAd6hl6OoSL/oEfh7Lm1jXEkXNAonmfzo9S79XUT
VtWC++EehPN3bk3Xx5RdHA+xOZr1SXCt1sXh3No40p0mqbo19q3tz/JgutLqJqQSQjeTKYgwtSZ5
2ZY08AU+Hfq309XLGBiXakn4PWoFz60wvAdae3td70m3Nme0GqAge3ZrhRqovt9wrV7OfmqZiiSD
8G2GddJOaoiNgf27bAOd543MZ2PaVdRuswJHzjZk07MmezyNubOITE5PolBmHSSs7pvB9ORS5rrz
Zgi3wFpQTH5lIntIFfkgSwX21j19jf/77jZnppegTYksx9DMHpMUUyu9YfKEHvNjX/JlWTkS/FjE
fz8vumkgWvBhPgbmSFqVmYdVVu10KHdMtd+54Rsfq79vOix523GaqLHUiaxfSXjgRF2SBCj0Vp2a
5vT0iIgeCyjiW/EN2keS0DzmjAKhHHByhJ93jTjFk/xAfMqr3LoON5qNIreANWynU7rNOXxiIkem
7IrqtVp1o7ga8f56D+d8T4crhLv6lGceERHwGQsSqfAfcilxtLK7Hw7GyuUvoe+268385sDLxEx0
Q/nypGMBXi3Fhv4L+Pr4QcqNWmDwC0SY1Z6eF+mJ8SW66qNb4HxsSzLH51J9WvZP4xiLlGJ1zen/
sQvOzdnz7iWquHJ6hpPRMIwrgLrLfbYDDEoUw43wJxxRxqdwhB/bRzsS98Y5e9VtPa1FqKMsA0N6
MgDMLe54ErOxtHYCCr0OyG5yxM5rAnKH1k7f4+58dmvQNlLh2FbjCOnBIHqHvDa4Gj8r+p0QlLvT
fpstTF+M26IkmN3N+o04zGCXy5hdhTSHVZqyG/rtYg4VfcMxW4X7KD68XOl+X6zxEs2uEqNb9I3R
HWQUZ/eClqBQFWKw4ypB5P/5aGYs0vjHqve70otUkl24ddPCPtQX4vEdiuHSHKbFg8wacugfybYz
2IyBzkrv7fzg/Ct/Q7oo09BSwkxSds7u3+MW9kjxDGEtLz/lElDYwfvRMqTuJUXPRBFTA/XwVI7D
hoMd2+8BtGx3o+OFXa5GKu631jNGk0OToTABSjtifXuzKrxmiroc0aIdh/RqZniLEHT/mda0YDpD
9XBQrdZcyh0z6bFu2Y5NshWXCjbc1/m75OUw/6CO3zF3aptmNdXndpfE06H7Gbg5fxDjc/JkJ+Tt
PZEaCkTR1URN6he6AlXO0NgOragattcCSqLLSJtf7+YvT3yHg2j1JSrFMmTeUXObr6f8XUbUgs9E
/Jtyn41HiXLw9gDwBqwp2SsyHDLvpYxj3iyVadbEnIX477SOQcc4FfuAwsp6yeQYp3ii2O22hcjJ
oKHP2+vxEf+OBekIlVjhVY9iMKHbiLcXHuZx0QJiXXp/R8dqwQkGVuAFmB+eFW+AbcX0gDY0weUD
9Su9IiMD4WalkQXpeUcaDyyti1ynwq8BWlRqF1UWUEMVxWLYJO+nbNRbxoHQeQe9bDZPCbvmOD+V
Y3ft4pFcv0pechwDBiR/cL5WTUxAzHDkS1eEjflIysWi3LrKvY0s+BFwzQA0NS6qdlLKXVdseKTd
51DjbAmi2L4PSWGjxVSkffWNs0tgQ0/0jLM6XvYZwlQbGSvXTuFyVLW8txFn4T/DR+0zpBv+a8d4
UGB8WLowMRY0CjcvF7WcN/EUxOWKE5AEyVvgL3crf6LrL0msYN2QNW/Kkpt5sTw3bCmJwMO0eA3t
oBTxX8znNefgLkXQ1gobqf3wx/8Zi5y9pxBUf8WpXFWvf5SJIzq6cSWmpjoJUHGB5l1LWckhrquh
kFyHSR30BJPAI3wT2EmjNlwYktd79MTvZ2ybcvsPw0QVXkx3ousPZKO8G10KApaFb98UlYC/UiZ2
wF3luIqwQkfr7ljoYG02R3lsJovGzwhPMdMxskSzdaB/Z9nI40SgSvVcKox+r33S5gKt+iuhT/fZ
hnecNLrk6rM6By8L/ZvLxXw9BC1X+OalAWJT48zPsq+eJpTX3kazBX2sfpH1BSyPBKryoNmSXwkJ
zWfGMgokOxZprtF8Ixw6BbjJlHvW9VKUbBatqEKaU7RvKTdfbc25MPtVYwGtkgV+wBHQg/dacTEl
7hbOx5EA1UTr0qy2MIMs9Hn7yiSKnzhHALMun9j3EJkGQiD9ZmaxPe4kt4k90eW8B0LcmvGVOfY3
vQq6Iq6arqs1SwEU0jDOaakuevl3gRDpuT+yku88CEghgVYcboPo9isw0gaUYbI6AVU9YUYmSukY
oeXJeKdaXdP9Lt1/jHkaz549pRzre2Kr9sMSjTgnFYX/0pO2UTvyRWQ8qKcxD9kmwkmUl74aSrlM
9RuP7WGYqWoEzwyPjsQaFeo46vg0+BCnFPCkC89o9JaBB3r/zkfg0Qf4FhZ05QN4VRg62qxK7kv9
R7SUKsrgqDS/Q6lY5CzkZZbh/wSOy1NnFOplUzMxsGH0wUuxmK3vUr2yOkr9prbgeGH3JBocqb02
EUiJN2Yg1tkT59ndUaqGaIzuEij7JTsJj1YcPcPpR+bYuWI5rBu1QI9VSPpWH3uVGzU0A/Bom1QB
kHmfr1M5Zpr7mvXArStGMnO9VTC0R4+YjxSzxv1/h0bRH3TDnB9ATTmrwVWQ4ujxfmfX8jUkizb9
YoRDbL4eImXwVz5TnlWuU83N0noOTGvSn76WcMzX9b9Mxky1liHp5/NeEaSIjoomA7QeWquo3gC/
+WoEgA7WhRRPrj4jGk6uvo/mkHgh538j0+bFEtojVZQLqNjuEmnmNCFvRPFkX1cQevbVs9w1mhPL
kfVovmw72lMVa4xA8W8WcXWL5q/D4ROcAT1H2oqEyLF1uRfUJoy/Vx0d7U2RWalwFznU4Kq5B27K
yZsvPjwZ+/81mPjp9WEHhLz3wmUZgRY/NJfT0+0k2dxeChzkty7aikKwiV0tULMk+O9fOAo7T0iP
ENoSdhN4XU6/Iu/QKObuKSJXDbDiBLe04zvgmRJv1SFo8NpD4RutJJVNQ+bgZFdvqgqWtv8PM3s9
4OWbsvoTJ7fe9S7JpLNf+DTrYSMMAC1elXmoEGy5kQOe6l5YYbFXdHYxa6ZSYDVM3dXMoNvP3lji
XxGIh6Sun53V/UjEvDcqsBTyrslMjIvHPFENL9ZCol8FMy0S/zji0IMb8t38O34u4kk0AgOUg8Ew
99r3VxBCnc/Q3+Foc4kj9ay8SfipL4OSSZZWMDCs7QLh6U6Kk3Kgw4m6NoWoPg7gxy+OAfXDpHfA
wXmFGZ+5IVywbM1Lc85cxVzRdeGhO4ZGmbvbB55G9QAsx5H8Cj9tcEToorTzQRxEHdYXW9xf91Lk
ICSxbCbZD/0AxHPT7xtvdGdoO1MoOmAFqZg1neGz+UzqfyjIm3OhrUZ+GzrP2uuvPWAC+7uiKmde
4WxDnf18eFyvNr+eCJxG8kcw8AkCa5TmJTMyQ1BUkeDf9yd8gex5cPUltEBUgsP60t31VPL351WT
WLRvxaxkpKZzVhamROMseR1dapU8jgQuxxX/SCaJH7raijturram7gVRWQAOcWY606U8nJI4oIaf
qzFL9cjNuCAIMe3lxuDsKXRUYIIOWe/Pkgl6AW6KahZsj3G5U/nrysXqE4T04GCc03CCkowNE0NO
qRnkfrY9FUSzyMVNUloG42bSFLNCSazdaOsXJj79FURv+emQAUrPiSwP+04ivze7GH4mJi8KiD47
hSVR6kEbmYRycKhxAiglQiFQ8bK4Ux3fIDzBmaCGozF0jgYhRenkqEbC/5jUXwS+X8I1SedcTerS
PBIUSqvRsYWjvMdMhp0NyH8zUT8pG2CC2EJ3FlAJfRCJFUF7YHo6tG1OWY2PXliQSR/RcDdjBHdN
B+qBKPlp9SQHMNaBxByEXa8zjutpDNYC+73x4mMeHVJU5+5/29LBdqHcBVLIx/Q3GnTc9Yn0cJ6N
nBsaPK2Q+byYbY1/oLBGPKQh4FCpr/HAI1qmgiyIXgEty6B64BqW09bgjHtRRm2dcUxRwcOjQ9qg
3wH4G6e1Uas6l0KX+c4HzhnQQMyiwsAE2vIIEt7ZeLlO54es56Ec/yIbrFxS6tNykR0OaPeikmND
5j1PSIKp1ABE5Cl+WLrZayrQQx5NovDNxO0AiIy0ZMiDbrTtOAElMpF9M1jYs7PeR4Wq4agEyPyb
7jBYCVeCDGmHoksBfbGhg/m6mwiuNSCvTp0vv2bc01BACDeDYTNlwZf1GUA/e84zXOB28HRP++z7
RkmIXCobfGx7UnmohvTPrRRSZ+o0b5FGhOE9fx+vnQo7raRYrNCO+DrN7a4GypgV48ZTAQ61oQ86
K/zR9jhIydyUEZtVFDm9i0rAgBMYqFZ4wiPfl4cgw/PvK2jRf+25zefbWSukxxUbE55xlwnjLa34
0ewQp8Hg8URj38OUK548gXSrCgR3LEedBUZx3LdNklpB+G/6FYfR6A+NZrrbj9zDgbY04aPNrXyi
yW4PByNX17TB1d8RMWQjkVhBOJwiC/sKXKu2GPmNMWxRK4sfRcnJqye9+df8Bg7qcNR7G0goIfrf
fx8YSQGRkqhsA3nhbfUySkT0chqyo1stasChGc6lziyrF3wzBMSZ1JvoAvYVeEaq0pjjbtg1VcBM
mKjrNWvonXk0oLDzI99jrXsFIU672Rvl8i59f5jQA1igK7I1n1KrCKnMBQiUkpeshtYfXAyrUa0Y
WCk/E3m+7P3cRTFqQDJPB3hPS7wnqDhvukdDQj+/HhzBR43vRKNQFAK/TdKK3eaXR3xVsiscka7Y
lUZ7w4VYNA6+dxflJyF1rBGPJKwQX5WmOlEq5vSSjnx4UINQiyHXmXwV02NbsiQaF2i9nsO8xjSd
StPvUiyvS9aCLseERrcncHzu33+Hy5G9lqHd9VMYqFjNrraY8oc8v+i/n6/I/IM00+HAGyflSyZ2
AfMaG4XzSmBke/lO7rqXu+xwpNaZgTf8eY4owCZ5i35nkH0HqtwT4HYZj9P1igCYocZ9VvkV9EXO
WgiaAz+1qhJ+HEeo/lMN9jmk26zu4pyt4aQWaQdLpbwONJuvDqA8B0BNMtJVPL75amqyAjoZ1/P/
8/tFEnjpNvJ82YbC7pbxqicdLZ0FwGLJOzUvKFou/CZC8JvReDzYO9V3OZ62IC+8VJAjFtRWet2j
ek+ZVCM+Aiue+YAnLTswlsuRp9Rhfs+q7I+l1p0LD6Xig5dE4J+AuBGlPjPctNDocp+Wd5vk1hzQ
w2L2aXOeJDmaIJJQqcZonTU5mXkO1d7Qz3FfeuLGuUweZsEFQhCbNAqcV7UROKDPz4cG0A5CS2NX
ymR5LMlXJBi/WehxtSgfZOZFkghkT4LVL9cz8q6ulQkaGl4s+ZV8+kzgL9HAPjKYU5WXASMIyUYU
d5gl6oFSvItlTJhqUKnePgRdCyWkAX0z8Vr2rD9oMUh3dUX64HU9bwuoFvMk/qPO3jxcZ1gMwVmj
S1w//QWCzCcWaKFhElsuCguiZU5uPabEDUYmnVpkotB25kBa4jqaUoXbOv0sCg2DKBU5jtzADNOv
QTuNQn4tZP62FvxbDwDHOshYXvYVQ9jGw4wz93dcyEpGPe4wyiTCkQeF9mv9PlId39EukR8VEtpQ
fC5tCMS2ywPUyE5fLf4XMoH2o/p+DuNGcRcDzhVKkxsik2nfK4wjZ3SqxcJkzmQdBu6qHLrg3EYv
876ApWtcLI55nr4cfMsrvptbMpI+uOhkvcOtwNWSPPfW/Eqc3shJeBUFH5WuOhZwV3qCGuzYoRCk
gMXCr2Geq1OdFBNJxHo2FPGwCeVx1TOs5qJVRo/x9PCj9wHg2qVq64XCHSIVTJIDGa3R/Yde9y6h
KyVslDQvtjcKkUa4tGJ8ZWTIyxNeY/1oquRFiYWS5yaZdChQA6P6cJgWowFn67hnm8Un1xYmpIeg
YtAKCB8XTnSPJnHHzJJI/KDgZrdfneW5TD9t3mdiGz376gNiY9LlBSLdoV0z3nNFfWkK+pIcAkgv
tpfVWUFd37dzYFY4VMxc3WcWwQbb7KEaFDwAe5Z3nwLQCqfgZRy0caYK/yToYr3qwIWhBRTClFkJ
rITq1I9NhnSHlyNbz6zs7gnRGcN1bYmOqEYtvvh8dQfVLh72z6QBldu+AKlUMfwChbtXI3/a0d+L
YNUpVA9T9WH5SOdbWdxHfOfO9SIKUG7QeLQT/xchdmduW8t8JeHeYP5AdS2rJdcF4JMPK4HxFBAl
71K1cfQ2gj+6CsLb9MaVQCEL5Lzk5CxmtHDz/V/jthCj7atx2wardIJPfRQM6f+2xh25ZDtHBX+O
Jr5DDt6LhQmuU9F8Mta5oAgdqaunvG5HeAsdiSvPwAUFEILEXvSHj40cjetBfaTXwwFpZKUVAQch
ZfyNUFoAtjxF6VcpWhRqCpqAdS7cupxVR6VkluMj4aqrEaw/1H2zs4md9jINTjuOVKqWQa5zW3wy
X+xIjmhxEHrX0i7vVXoW47sqxCcXrxzZnItIp55khRoAryjY3Zfc41rsCVn8TqDGVfI/xHGX6QlD
YhqgY9KCCicZOh67XCKGKho1+Lr/vzPDYNsw80y27BDZYxoCMFPEK7p7gWvtr3fxq9BSZ4EL77jv
DfPCr5xvoQCNSbHDTY5kMCr1lJb2GDsqdVQPDFzNeNFIi3EiutDOi80YV7X/+dAPCzquiCrgLpbs
himPEsZtm7X++vHDvMecm+Mmy5gpKl4a6uGcw7vLIPrGq2K3XGYa86JjMCROLabTJudL26yd2Eid
mrbmOi0zJMqVWh2E7TGMRA7UPV+FMQrvH6CXnQNMZ4B0lSL6ro5TtdWwBcUyBVAJug7nx6wyos1J
G6rAohTJcI1+ydJygknKekbHbyhqXfz7H6m3jekxDY/YEiwff9qMxMGat6vgvWwJLn7QfQt9bEUC
Kwm10byCnODkmUjU5HKQRAtD4doobmjarQR5gsplH80MwvQqcKm5r1QegRiOny0iejwYdJhoXW8w
fey4Vf92aeyqosjXn8un1gWEu1Jz0Ck/827kpfYPNWX66LaNfbjgE7wXJu0CGHlAZ4I7Kl3782h+
drAS6MT5Rs7jJpsaow6zDVX+flhyo1C3FBsBM/fgrh9rImfIKSuyUPXcRRFKcC6jIJ7uqiE6oJQR
CgO2iF7T46aCJ5uxgTdRXkrAKWDohh7be7iCTmbOs56CcHGB3R2wg27TdmgM/jETmpxmuB1b8MYA
hB4QXx1IVsSVtp/ZaoY4564Y6daiXPdkQYxujQtrufnsdx3dMNIaQ101PVkeFsvS0cPcLNtlCTJW
yzUoXr/ZYoUxx7VM9ek6IQ74oR1yu+daw2Kxv1Odkcprg2sjThHOEe7L0f9bLsfNY0SDv/reDhlx
7BE+iA5EOHPH/WMKUgPC90HDgz0IWxMBYnd1DkoPAYsMH4ha9bHUVXKgAYoWCkQIUVwRyfln7HCp
kB6gLcb0ZY35TkKkxl7j7W6f4FW3ddx8Ub6YdxOOz6PvtI1Dh9ck3CN6ylb+Dg7rAjzJM5IOkIb+
syzRU8iA7CzEezIXRQsF8u6d4sg1r8qxEj339whUECfsqdmZ9vmZtTzgTGbpLFn4naJ44eTvC+Jh
Shs61a3U3cxMpK0Yj/wob7kcS9VwiezegMhb1wnwXgyIyVmDYi8x9KIBgv3WZMdiaTA2giX3b0l6
V4KytxZte9/kdzDiyvzevw4ViheZa1wno8yRjMfaWQStuJuBJFh3T15Von7GDhb1rxyOyRJ+xGPc
QH50EaLSQjvZepgvJwDFlBTVL6tmyueWIeJwKO0cAVlnETKBlh+wqAAwzVWaGWJaaQSThfNzepVw
r13nDi0ICiNF/jZOxf9XqAVchCJwMLM8lhXtz2MoCdRnyadHHg5RSd+dwpsQ9jVuBVUHLRd69KcG
/kzACx+hHHJXpahfa4nS5TMHaM1325ulxoUEvWDJKPtC6dhvZuzDQdy7ATSGZdSypOQLcohgJKjY
P+oIWTgG4tzn3yEa+yUJfpTIyS/MB/T+n6wFr0iQ8Mr7qMb9lbFZ74Vbj7twQEHwxfKCreG7fMv4
XM3O2wdW1Fgz/stMn9NmzJFRl2o8pu0BTxtFlo6iT3aghEq7yRA+bdG0lznxQOEpuzc6p7lIwIQ/
OxQQZQ6z4CYc1SfCrh9JI+FPRe76QB8cBcump1N3XVek4qgfNPmqBv7tBXeIZloEKCGZipEcWkCB
sHFsqEtlgbr4seUpwtIb53QXzeCHSL5BKEyUWbOYG6hpTGfoXzjxnDxoXCqDw3EG4TCLKSQ6L/lj
/VLlmk+MaZhkgdxkx5+DwvwnJqOBlZLovO0EyvIUYRMUIiQaQYmkm1MowicD2/Xb4UOIu7zzJeC5
P4mUJna+lz/Atng+OqEfvp1/iUc5Nc5JsMeEx/6sgYXa/mP0WcvO+Jv1TiMw/cpVu4DYiY10numT
2d0toYoZtlziJSrffgcX3JE+SfI7ANUbAo5fuVVuZdt2pzU097mjOJ2zW7yRAXCZfNvuCJSfh5d0
Y2bz83I5j+459hSTpdip9PZtoQ2L1ec0fMnUoYr17EhiayxvEFOirhXvt2iHFtqkIdinGxFRku6f
hWvTpbHLc5hm7WJXL0tyX81gMFgAk9FHRSAExpWyxxUUQlKE/ni5Y9FI3+gfWitjNlTdQVrCZvFP
/QVxBK6R0he47ONfh3ywG5cc7gKgA59Jijw+FZLvynaBOAzQJl1SukV2pdFUjJzoaomMGOtDu2gv
RRY8k5d25j9b2rBlgUX0UMyVpbxtYWCnvPUQueUUe29u+tOhtkylXDSyrnFoxwcaCZ/RPxy3oqkZ
R6pJ57quNJuUP1js6537ZbcE3O40UEws7CiGCIKSn58v3hGUVinNTW7WbKggLU0OU2M+MDREpAzB
tZMIVkodKd89/lqkLwLgjZaS1YH9IfKtzngwopsop6yGRzYmNnj5ToTYdF0xRxq+yNCRCxq/r9kd
R8jZVcH0Eguu6Uybwyylw2JZbg1r7z8Op0UKMaUxnXi1HGfujkfX/weJh6nWTNDy5wcJJlYv3xG9
pjoxC6G7aBro+lGSyaYMN9QK+hGf1q377oo+LbPqUB+83AnehP8777EhjJxLbB9iNm5WICkjWfK6
fWezIja52KQh6Ci5LD/W0dFonyYAWPytDhzdzUWhRKa3PzQ5JwwDiDrZP+sDn9ZRsteCSCZ6Q2hj
Yoo4nLLfF5AmUwoNfoPZDYsfWyce3km0xI/klX367J/q6CFvjQ1DVetgxSRhJY/irPAw7kuvW/eH
CVvN+/Ekb3+lYmnLcHKCGpx9ci4gUGZ6q+abQowuXFH2TeHfEnT1JQIGbvAueRbt16ZNyZwWanUd
HT82vbciBIl1HzDDIxloCuA/SlxKSEQdRJzeRi9h0EMGzxqhPBXMs7i8HCo8LpEg3RsRjIGW0wcD
2x2M6oZps9FZlFMonwAUEp+TgvjYJo8SdA+WSsC4AOqmF1Y7ftsSCU4SjkGyVBQY8nuvcp22LsWl
XvgIah8XnV6l5NHD9PbRZYERozMNW1uLhRe00Txy+XqLY6hkLAz4vrgE12Y/3jQFc+BjWPZ+cmx4
4el4xJIQyCulOQnihojXxbcaCJLv4BX2E5baP1MefNoO+qD+w97an+T5Unr24SVpsEub4zugeSED
QMrsN5rOFFSJNig+zlInSA5n7X99TZC5w6mDzssdeEqRKkumErL+0z0bpzjDaYcE7Y13CvWuRJ+d
4JXfhhjNFQqH0EuDqQJTIYvp/htVmkTugqloqCDGNNmiLmcEuq2ROs7M/RtP3ph16T1OhMrKEaXW
srGlRU5/3KSyNa3Ds8ZxFp2ssh55MNa08+VpyTGdXTxaeoLJUFXqIkGn9cKqYu3HLqU+8KD76NxM
kgL3pm1lGByk1KH4a1e5jzqp9gMJlwiIwnYdv3Famxt6LAlujQyJIX8te6cySzwdH+eAE6KZXh/Z
MuXqvCAQIYfwnwPMd5cEGib6xiLMDB1IRlt7I90Svx41n7h6s/I9hZYRGH0NsEtAcVqAmy1EA3qB
cwj61NldcvYO8x0+uWpd2bB70NVJa1ogrV3AG23ObmXmjJELEkkDpO8ywLcjsV3VTEuq2OcS5BBH
Wy41WLEX1ehJRCGpfBYIj9df4+qtuFCJsP62KkAQGzRGaTyIrbw/1aSTuiKyGcQjl02TUfz6maUa
cwIF1/14YL4ZB3rkPYFrHjn+lEcGCDstbdUCaVgiJ2CHNZax6yhaLordx24UfIq+2rWmiM+upTG5
Ve25KonnOW30OOjb7zpr9WHtNXW5j4oB8Qw8ejfPwXwrAOEurQdZlj8GjZUyegEIMKjYvbQBirhQ
Bqx4TuG3xpWT9+TaK5ZQJBwKqJnxkZT5fa2qerfbkfNakKwWIuUmUqMxxCh/Ju7olXmryvvN0mXK
jqTXf/YIA6Q3WgPp90hTTJYXjRRGao5AovAkFq/AJRjeV05zIqRxS/brYrS6K7qIwMiK6g3iHrl0
FBL8CAcs9FEwZrORWWgFynENWAHt4IajPvHSLViquydgcbxOlDbXx4f1HkvtWbA04c9/WIa3fGXG
68lnHQk/jRN4Hd7erc0oXSFZYtJOM67OWTJ8r4RMuPqH0sS/lsUtH6DOnskqaN01xFje/pU4Rlrh
vAPzekPdUppnWH5BI5SI6cJkhZzhbWubZ6pI7hOl5AMxiyDy389SeiSFd5Vhb8kySV0FpjTscLfl
SCMFfGZENaolyHXii13DYRVJWLwbsPvMIIgLvMVTKUVQr4KlWsOnhszQRvqgybiETje6lycEhVOB
zW6m6P5oQIuo3ncEuh4DYo7kaz8jqR7FSQoE0vofA6ojIRa6uKxoBV7a+/mH11/NxtuALUxuXUc3
7TC0DhsSt9oHaTp5abf+L+kiAnSCQUtJU8Aqo13fDf4fulcq6AA1mCJ7GzcmeEDNeOJHaClHswev
yj4AtM7wuEsOgqZ29McmH4yVL18v8D2U9XUXuqXlynxiP1Av8TqH6ZBVTRHj+2AZ39khYjKU5hJs
Sxwtc9/GE0CvjO8y5k4h6v4Q2jYKIbIl1Td6O8ORB7JgBI71vuVk1LmCyN1QirUVCyhtKWxDznY6
dE7DtrOg8TMvZaTtU6HnHQQ97pJkTY3Dj0Ubt9Vj/rC91L1FLDpXpbWVmJT5GDxMXd13rZo0XF7L
J146aKM/kg9x2qp3+TeS5SyYvypFEpAXUCJJ9Tsa/pGYtc8MMD/4fXp7nNOQrpA/AXx0c6BpNcn4
dD9WjeWmnm6rlRHVX89mD2KhcVbX/qRxG271BgfyykeFwjiVxVwv7fvheqRAXkRgHpzRAMC2F1Go
ABqyOAfrTecTb4JOQ6TR72X7sZ2UVsvkDrVp9tz1ZI6yNbixlgd+osU24xyDXwp6idwZiuossv+I
3DL12EXfIvxm06ki6davjepDnMUaHiMCJscWy9qj5d27Q8kwaXIHC9TvMy7QfVAFbR+bKEsvIZZE
JsVl/16Ix88qa1Hf0fQqcCh5uzgt5CapA0d4PAWxuahWQ+6C0f0Kkb/Bd2I/gOIYVlvr4V7cfQzg
1WUxoGoR1nuti3GTLVGE43IGLEXuUPe/jj9O0wb2QYyZLvq/8wNZN0yoIoG6X6lAVRgZ/Cmzie6j
xTUq4esWSpLGrSd3t4WOJqJK/EBst0oa/t1CzWqU+oD8CnaG3IWOb0Gq1XBneG8sA40NDIde8Qo6
ZrT7Hckvjq2Ai5pRdm6lLQFbtNKlRm3sjGc/0VZF3wzLGscnPy2sZQTV8WB+/E9/u/4Dr1Z4qRlv
9zg+VcSd5CDVqP18Z60Eyj4V8dPqe5dS/+CAtWmcrXRgBmcPUjuSnesCa1vSLiAA+1rtnAl/qUxs
JZsK6Dp0XlzWSC/QKWJn5wg+YWKxQMRobDiQhawhyeeVk71cw3q1JlmDAJQPBKOpxnaiZKRlHWBt
yMIkbetkWWk09URxwvh6NSFDRW9wGU0+SMyF61N16DukGE0Hhh6lVaXuqjXlO2Ppfy7E4B2qhaHG
pi4YW6+fLBOB/yr7vsi6DlzimTYPBvzTZMiGTG+nohU/RUlwLOMuYIqpFw6Pf3dRAJW1xT59G2dm
mUuxg1kqu/AXfXLdgeuYAZUzkw47ipPvDRRAKZOoteyIsQ+53YdoWjAKWLwviAr+q0Csu2KTCBrY
0X3aw8j4NMoHHw6MOKzTbjSxggNyy0LhdQLoLuygRWIYSahxkA6iSJHD10xJfR9suaDTSk1F5zh6
+xt/UTy17S/rhw/ba6lkXrG5BxfmtjYIA8ctL2dibCWW6e36eByAD+pDKk9bHHD6DoZfvN/N7Qio
vAPNpOsONEmPHmeEFe3gDtAgW/glq6gE76pNb70Xr07ePvjWcYCHKY68LhKbzOuvuRz0I6HGNXUy
vR38UPaSK38QgLI0sCnpW15vv1yNiPt9+nj5grFs2vnR6lpaBleM5/oR+Srj0Ym5RAYGb6JRh/rp
YiyYdg69JEjJQlUiGrxGC5wV/TmwvEhROyWKBGQBW9xf1+Pt/rrbXvWkKIcMyyPRp59gSEqqor6q
WsZei6FiAS3I9eAO4Ie6ChaZoGAwxGAe8LwFdOEd3Fer2APCfBFNwEgeQfz89P2/HKywwLKRfliC
L2m/65L8rEghaY/Tbbd7d7Xbi0kTlYK4bUWGKatDuv5oLEqkGDfxHfTXsu4yDcWB+pkz0YtiWPZu
8MlT+Tv3nHEKt8o/aId/00mnf62Wo0+cB5GBbgCGaLIelBh3870T/zZnaqXQWtPRLTZlhxd4I2gl
gR9he6za60YHj+6dZ7Ht+aMwIZaqCtaowyYSHbfGVay64KUvzlSqX5rMwkKeOXLU4yDWevJa8yGe
MbsC6d2xeFDx7+HEiNaHuxgWY4et6URJaXE+M6b8xXw/uDtodAVOoY9d5/f+W7fGa0h6qkkmEzzT
sNrXSyL7Vf40LsbHxbRHd7tF2i4h5mfzKB6Vt/gGNOiD+6e5flxH/nqoqI5StwADmTAdh31MU1/Y
UtSaUCwzgOvty8KlK68QvqclD4Lt9NZVYoX1zvHVTtHpG35XRz7Io/qWfU7NLaWP3kUrftwNadXQ
eSVVYey7BaNGViffJ03mT0GbO5zjC14Sk+AUowvf/NFXTnySyvDR8/0F3MIx0eWP4SGURRjW+wOK
xUfkLvV3p/0u1qWEZOZF8WtC89X+jVlQaJpo0/bHgSHy4Tny140s+MkJ3+CkV5G89VIcAJedBJig
pHUkiXqlENP/UNK+1VPh/UjiPaN3Ct86FwBD/WNFh/Y35edlnJgik4nELYALUnLEoa6997g9fAtd
jY92MMDIltVS/Mw2F4Mmo+e0s1X8P9Vr9sGbHK8GT3U5Fp7JnKOgA4/IkfjIlwX8PCR2s5k1aiXW
3w486Maml4hddCMPtn5RZ+e+c+FyUDqW8UsQOWF1rxJgep+KIPZmtWTOdR1m/WnL8fo/VW3zFhuv
AoE9pD6F71l5QExn7ijmQO909g2SLUUCGDIkhH6lc6qwgHQfMvGIiNST5elD4Q6CEMfMTf/gQZZ4
EvJdHlVvf+hdC2yHZ52yg21PqGPUkHfFssZY1VvAVsWlIfnp5rwa+vduyPownC3dy+0GH9gI4icb
/10udxmRTRJiwP164NwkXtvpx+8sRIcYmsnvEB576YEOJpydkfNUrmAVSbIbWwt2UNVHFqbO50i5
DbmAG6UMC7X77IRh5Qm5dVqHwU8ItFn64S8CtlUAlzXvd94cH0t9kXK/g+rRAxIzs5zXk1bxm/+O
uRd2pv0CmwPDi7Fva4Ny8SjwUyqvh+64V7mNlSQoF/2G5XY27sBLVY/8aMuSdHujf8O+hdTXLA4n
O80TtMqTwDAOil0s3kS0M5PtLMTxya20P+BQ/7UfpBkbZDsVlCOYjkAr8LTbyBVfTcknm7/ht6n7
mFzlQ+MreJHiAWwAreHs3xVAr01d08df0BptVrONZDZSoA6huj1qOfB1ZMgQsUb9Qc1sD9SiyLWy
4R6BNbWtEouEKMtcBm6qePf4Kc5OUyax/+ewTbyU3VfaeClxrK/C1nWJIfoRtry6OymrwTaNoHEF
RTzYy0boCLo21N+Ag68iURVDuZ2VInnn2twVUJJQHAIZvbdQiliRC+pYhkFu2n1AbH8NUNydsK+r
mCkQkdIvh/qTOI7c5DaTkElUbY5T620+adTmDNYJQqdxb7VYkIFfdhpkKhFN76tCmIfCdc9/0tL8
+gJ36b+ssjdDf6Vb2CiZkjkb/42LZSyd/4/6Yh/946lZs65ra4MWDMLQW+3T7GKFqRMw1UUAZGQL
5jOwCpSvoGkar4Swq4DYFrtL7wZKxyMXzmsR3aD0sfGU9L8lmeQ1ht4e7IlFZUSzYV02CF2zHICn
Zq0nDhbxb+UzIZVXg8cuuEw5z0tgT+9qY7PjZUH7xM1j2cBpQDVV7yqjKGSuyhia21tw6sqP+XiS
qjzOnywgmmkWWjmTYULknbGz0cRwZW22yn3ku/B9hkiwV677WVfuPbQd1+ZQl3+Mq9nC94jy89fE
qzWtMl+aBhfKkzA1ryQO/7Vn9Q7vfFkdJr8XB8BxyLZNh73F7Y0bwZ0iLLDo1e1cvPuVkYoR8hSx
UeDCcyyCBYHpbLlN1yWTMLm76BPVI1QP4NDvFaDQBe3467w2U7E5xShhOry6cfmWxhjyY+CwH+x2
rS4vwGjIEuqFK9UnloIy51E07eX1BlAX/idOwevwQZKxL187M0so0UylM0649ZLKKpVgg5DWBYCr
ig3BGIpr4/132MRg9fW/hR92cn49xOKiHB6gEo3hd6te3EZ8krXhW/KnPCnBcpZcjZxUeApMMHhU
EFZOq0ttdmpH4xr0X6wEleHRorXoCsZj6zCQtQ6b4lfO8lcAHii20lo7pkHRdbKzDqZe1KAN+r9w
h0ipfw6eB6Emd4ED/5OkZnyV656dUQW8cPxEohMcjzz6WYBRg8S8wubWTeJV8IYlKVJcdkDx7864
+Sh9MRES26xr2+zvqz/zrGkjo1SOPRrGeZuHxPTLrkjF8Iai6lz6jM7LPB97DeS1GRJnKMhn3Cde
ztoAxbOctKJClEbMpaaE5gvcErsE6qymGgrBXU2hEEhYcZu5aDdBPI+mUq7ITpRKNPLUt6Ug096u
8XiPJDrLzu6yRE0X1gQPjyI/F/E7nS7sISftce+cOCzQMT9Fdp6+j+Gp2kbqMvpMFGKcelPjm0NF
a2J70NuwYPUAncPjhlaNU2D9AwrNWq4SVu3pL1nnYa0fiGMyFrdushfS2MJ6d1AtjqtgHjLYP2+U
n4ONnrx005n9T4zjbbe4+LxYfO0l9Ss+csIxpsr4sKAzXbA+66G9ctFlkobzE4ZIfXX7QKpEIqwI
EAwIuvNHDj5+fEISKQdcEouGboVJf2WlpunJ1uu6iVu6foXjpLSxuIIxKptc4RtndCTTsYdHwaoS
RUFREIL+UUVQPG503FyM58jp15HGFYWijMEZanGK858JsmC65ZbBiztFtN5coAPDJMJd0DhTmPB0
JLYKY8fslVIXuFdQqDtZAJtNHmPgxC3M3zugL1HTApinFxeXD9239qcIXbqD7qmjjsSEPhmVCSsL
tEEwLtIzIocawV3cEo+lX0/LCWeoGdtbzqfPiOZRJ1sULujkAGXpjdxIjPJoclwnuA5n5xMh9rYe
csZP2eCOwr0lQScwrYygQlMJWCw61Xx+6sOWB8ycaRkOlQUmssNNnpP7D0GeWYMY7NpBnrnkMBKB
egNSxoH7VRqBqom2H2aTw6R9LqPyUlzbPZhmULRMbKKjcVW+EjkQcW7JpgGbyGC/ZZEy0HyGQIsC
LAgBYdcfv25efiCHYV91iy4P2g/zgqDtARQgAiPPMGmi2mn6+tDTI3E27rOE+4MYclkPnCqJ75kK
Grjw/Ne3D/kvO6YR90UujXOEfqbxKH9RIezghZ97ZCfFMLuK0YWu50lVxcgheRVWab6LO7pQ0lGA
jt1fxmXfRBb62/3On94MKGasWu0giS7a8gMNO1+kWPENGo8NPOGFsDs3+/7HQLZupwCtRjce/46g
DS2e2Ih7YnxUKu5t99QSfu0fOAOb22WVkTxnpwA3cjOkj7CB4SxnNBCI9G/AOx6ofQiaYIxDxdGZ
5zvxTfToBnNfuFBdvZZiDQZjcoo6GrXFEC+ZquG/7CMV/oNRCuGV9sf46zZuuQxrEef+QYpcCwKZ
2EOUtsnTH4GylMeWfMwZKfANH/9bLrh9AMJl/GsXIboYva9WG6GgntPpmopB5NBKy68+PzLl8SFe
PPN8ZBe/fPfJS60g55Ejysuu+brjQcgoTAk1H6UfluAHxibuMzZaGgm3nfoQ959SRrXKe7RfLERR
iAMRDbPW9AEbmZSeELCerctVbsWozGnRAarojT3Verq1V+gNgZZIqjDRIJ9xDhqAPQP26lgBk1dF
0pAcDNewZmX/0xt9xY157pz6Su1pNA0hnxrL6Yv9/O3QTZRfAxngCWgJWR9AbKshP51qW5AhCvn1
yqrFbQcOQpvFMCSwdlKeF/l+241bcdYEIZSAMJdE8xm8K/2wSj7WxkV3veITII1YzjvUoayaP2Zl
5nn6yuGeNMbGJ/sFUUOhP2Nf9+I3Gn89w0Wyj7Hh5D3m1fT5kziOyeGEMO3XGpZHhF44YKZK0ABI
k16F3bvHhdC3tzGUu3hWwDAglosW9VZbDYKd+fD/3z3jdfFW++a3YRvbpc3J7qUkAg9QL10GFwv8
Hp6swny16/4mxjsBljMOh91rsr5ibibN3yTZ9YflP5dorEUkjvzu15sIdbpXV4ceZmjPajelqLGD
S+PRzJTfJCMKYHKgUaKn4Yf8XrIX08SHWe0rruBtGS4xTe2qGK/MA4TThIB3JpfRRLIOmgQJ30a2
490exSAX3gmyKbP3cwGWdHSHZOwayS63euz9LfqIGSQOPU2v7W4aEEkK/3NQpzlZqn8y2++w80/F
tW55pKS6giPVTmqDRpn8DlX6DPtgtbsAG++iBn2IG1Kcffz/OCPAzj1eqyHflI6l5oZBZE83Fom/
x5JsMnkT9vgtJg6uJ/unfXVsV99xEdM/xl3uUD2beX7Dhom2uzbXTzr3TZsk73npBHyErWzcH4rz
bSHG1hNwiuYI1cuvh8llzdUZRLLh7GNatGr2LUY+/BXObbS/X8p7/gsO4JuFX0Gs/je0FJdJUxZO
ewrOQKbq9GXsxZyVqhmyL3QauV1Wq0FByFhKMEr6Ww0g7Baq9clExdOh7DEfZk3L5oaDy83GN4Po
Yp+qEwKCn5b8Wb3GZjpQYQfQ4yBzXNfsUqbmsacu6dueFlbgGWCGglzMbaSyz8+3s+MeU463HoiM
/ZA2ifyuSW8hySDdtbzhwjgeOnOPF32zU/5rvpdEWzXCN5dv4g7n8vRCdTpjw9se0JcsrEw5fvnS
lWhWwnuuw21Y7MjhSm3lufVMkfwHBVHCQwzJcTGx8vfF5dQv3w761H7oVwalw1WQKx3MiN5ozgsX
Hzpa0fFw5gb9pWnBep31R+eN38wtfWI0RzhRX0dFrboRBr+DwnGv+WW7Xu8KL2irLnEpbTgpiOC3
sLwbiit7cK9SiF8d3UPRMscx65s73nu6LS+bOVO0dpWjZ3OVT5jt8xTFeM6BLNcl1zVx4UPbdtAx
tDlTX0G9bj2oo02wltigp84Ta7dy17a9jdKmeHCKspvq8c05qg5pZvOlD1op1zE4W4IB16AQrbqH
yY8sHjTP9F/8OtBX8ng14efkRwJG3M986QXWO1nvDucbIOIMZo4Thdj0nEktzmMKzbnyIP4uwGeg
4sRknnZsi0iNP0KjD2CdJW/GMynuI3skCKHCoLH306KQ6x+NpCCilm62y9d19apmLvbkLRoRjfRS
K5oEyChfLbRiByLfxfsN/qLDQX3d6hxfxmQ3EDQBXVbHe6nEm+xVIh2TL2qNZkEFL47eUAwCEPQN
d4X9uhCY04NzAbYAJbzB4k3b0XwxN6JxMxqgeYuU553G8tb4JINWaXmZTpPxnrbZR9YhxMHXfoVZ
PHxOAEnvY9773YpDevs0SAMNRVHcoq4JNwuK5rXJXVP2ZeR5s4f67G5pj4j/jVlCt5xtUF/UbaUp
c4DADLZ4Fyp6X46SipebOGcv+Cnh0gAdCK3NGAL+LSox2vBLuezDE5YXKykD/Xd/GiKmgz0XB+xM
rAT0cH9LRHmPxtaeIGzwM1XYpd1zAo4QpoRzEh7mtmxQ3f88eL9jey1djALybuKJyjusi5TzCR85
0VvxQE1O/XFl/x8OmdqWP5amPyrR3ReZvxQSoJJms1MoLQQSl5xWdgsM6cr+/hgx/vMhZbNbHv1d
85CIHXwMvGL7XJ9djMb2bMJ1Xcky+u1WR7XM0pbpHHudTGZYJ0fOiHfeDMuEwn2D26QHgI14ll/f
AsXvgqWEzG6G2alYA1K/9tTfrVuLTbpHyNwJ6hnD0eiODjP5sQVF2IDVXMBZP1jP7Dchj948CQnZ
JCAjsKZALUmNpzbbb1kdlcfN5tjFCfw8P+auS8tRkVsD/KWUy7xtglnh9/vGNocthmDmC7ejNZjh
Z9CM4QFqpzV64Q0RkvMvqvHOixw2JjPXeoqWbJhbx7JkGk59Gh+okHkSsJxJGkf8OeZIFcbgATAV
YD3MUxiW3N8vMk65H3uLfQo34fTSvY0eYG6WdMuEd3dEeQw91eXRWaT82o/GcNIHHoszp/43yC35
OYxcGA6kAPvkMugwoI/CIwGbnhQaihYoOW9S7kbBL9WdhwymQYvKMZLMrRAsMveqtWZsN4EJzVfn
kDXtpk8FzzHkIMTlHYJciA+YGPlgJncbLrNIvhMvSxueP1e4WIiGBR1Ym2ZQjdzZVDThhjALcBJ/
LiPAHBzKoQxg4C81b3iPEZwOSpJI/ibe3724SUnV1j2NwiwSQYK8xG3zQwuy9IE99EzMXTHo6UCg
hMjmgw2LaiXSmI2NLVRNSKp5sGKRnue8N1FUJ97mTAWyJFkbulLims+nE3dGYy137VWxbZm/KNkH
w77GkDamjZh928vIV188381DYu4aSSi/DmyUlP+1NYycFtkaoWwExgYrANHSSuawDcQ8v7U9AtUu
TT7D5K0Xmuzfg9NXI/f9lkph3m946B/nMql3FRa/4kVf9LPz3YAc6mwctRPwMcRUJDKgLEi9AiFR
N4ucZ3EvUCH2tps/ttOqKqN5tzvc88tI9RJBlPbaBer3yB+QUmaxr8Tas4I5M+4fDWjxtyJ8lz86
s6Y/NLWWt4MfiL1JC2PfGpkePxu4ebVqENquTM5v5i/rYJJEJGkUTDM+dVk/FDYEILzc1B5zSLJ6
kxQLdWsruyz8h0aPSrglN4omNJhwDIvHU84MOtjhoxX0MMimOEZOAJNS1GFtSAFZ9UVVhA55AOrM
03QPvzT90xtk20SjXDWEamKYC33SnKpYHZTZKZT6P3sn16x/zqZdy0bKFUgUoBRshKRHfewWZyQN
Mm2JOn0tzpeiTZ0eQ27PgiqOL7DwKitGDqifhYCtgi9p1ciGUtSPNhpdfE8yHPFlBmXpOkIHTuTQ
/uh9Jx+/pciDHzQL3smHGpEczkp+xakLPmMMzC4AM77ItdCVXX+882W7Lm/bKbbCZjv0N33vGXqK
7VXmJtQOALuTx+lmYbUmTkQOgcNPkCJF1JCj7CIBRE4TZu9FBzEGp/HSmGNX28Tvq7CcVexub76J
PU8NXpxWbuMpkB586LPTaMWzsWr2Ix0IaLgDgDjXmapDXBIivi4bZWF1teWTNgQPbZ8g8vx/IlyL
A0ftevTnr9ixfEZ39Z4agp3yyuVUViulUKJ9bGiNFyIu5ip5h2mduHPHmzMwVn4NJMOTidgbom44
iNQNfW3gWBEIIu3sNSfQDye/i0yNDk0VcoBevm1RAjDjvZbm39mUTYF4Qp1zmfDkzmiBcM4oi9l7
ATlmByW3ZmmXnsPhCkln5hD/brafRU8OhEJC3glZfO9h0K7OijP/ykaoBhdMFeAp6baYEm1qrDsm
M0ft6EwVBWvgAPhcrjri41RGdoHwNbyhBn+MWh24uCcOzRKRBXyVEFlJHAmRJUWfGoTLGD50FANE
dN0beyITtf0UZ2LSVU2MpW7j7Rlah3AwV4IyvQnOciPtyGbxYxqx/RG3IJrfKdmhGl8PSPjzCESc
e8n2GiYZDke80MDizGuhfORv7V8Qoqv9Zw2/NR2EmqLVTZCvb73q0XyZRO1yOUnt7YJ9G4+Axo3H
vaVEQ26r6PzjzpLnsbrM2oSW6Gi6JCVrkdeL6K5b3IhHxm7+RTe9XJLy8QIkgx0QKlRT4x7vkhV4
lbXsiGdUe4MycUJlFNR+XXGJS95EjHiPJHrruiFznjCC58PQVhoFBdz4bjB0zE/va6tS3ZZfrMtb
v8QcICS6E5vWESYguhBUuW8UyzUN6ct1QNzfFX2X82yWfeCz+63eZJyMjwzQiB6l/XUgPzp7kFFM
8nW8fg4JbFlF94AH2ol+TYjZoc/owWyQcEY2XGZNHjAvmWxUk1pV2f1MczzCuoW37jHiULKyqqHj
bpcykQwa7Pn5qViWl+pRIQaOY2I2e3Q7bNQ4Bi3rK4Y4rPWw/c5FHCESstZFyuKE/C5ZInwqDXsM
fdMIxJklMIz8CLmlvClJFVwmGZxfif3QKQN22pl6N0oP9EJDFjcRb4629LJeTsKjH6ppdlhFbFrh
d3auB++LaZpFxHPw4dQEtudx94BNMgnFR1J28fZWV1hqw2ChKi9+YHIIAQUVirK+qD0Dxir36RYe
mk8Lt9WKASNEWMrocKdMOemd8Z3K29kyb09tWGMb7xQcVzq9WkvWZOKPuLjQH7UQsS46zRTESALF
b5BqNT7pfMfJVBeEmQ4iAm/JTCIHqQ3V9UzSjNRCzzdl0HTzeMZQxNmT57mUMpAwvWQXwOs+GFW4
U3DpaSzmbVdRbRKXr7tP/jd32as66GZb1QbgC885JNL4dWu52kgz6jMCpGkEt2krbLvTpWTOgHJS
anV78a4fBs+lKGlyPCo3qBel+u0nU5oMEZf/MgAlFhC1VAaCHI9qEDJfu8Cgm0Sskv94rQq4cznS
9zdBsrw9EQlk8Fk6hXKfDO8UIYogqxiwtMeeOjDvFZoNIfiOBbROwgxLYYJ+na88k0S4kbOpAIrC
whWReShO8zHQmb9zOfANJbote+cuZwGLmS5wV1Xs04vRBU9nPuZbeCRPoFtyhey5cNTBCs0n39Gu
H/NafZaCYV73VXq+sOs8We+6KTU7m7BWqW2WFLO4EWdcKVOmOwV9YYS4tFpvKqDq390ah/hKXZSF
RBNtdRVQHywtLBwp9o20zjneLtJlcD/pP4Mw4NCVH2hoTwG8BifPVBQPtHCK9jjJFRALAvphzklX
tpmonxfc6DjL3opuafcXMWxQWTFbR100yPkNmMLU61GRfjdehLy3b+Tx1Pd60GfZXL0pn3X4blC1
TNAy0F8G/bivcpB/FIZdKI3qmakAdN81WkFZf9pQmu9Afnwk4d8zfMalnWH+QzDkvOzYr8T9SNcb
7d1wkQwuT8udJSZ2eX6pfxmcHIAnNdabcs+XUvOAPeRUxkw4ByHaCP+1r0VKsgE3jOvDHi9nAKf+
hmG7L0f3W+zAAbfkHZo3CeN34Yb3q8ehhiQKm+Rj3ugeJPKioNOnCExO+k1mp/NeieaRgDT3B4Ia
h4c66wdiWByzSbEFmc3zQXbHVQ+doJFIAqZxuIR0uw1LY3tDXrNixQqdH9e5yDlaxJ4WR6UwvoA9
7+SGaY/dOSQVdzQs7M5MosNdtm9EdA635/m4BsM0bev2toyxw5YSq2/CTpJr/rWPRDuD98Ahttdk
SiSOk3DrIXIK0jyQlFICBrmLGdyavSJfU2EIIotXhvtTPtLSjj9nxyszGRN6VMmPBggUEhiWh9pR
ytPT1RmZ2j5QktRoAT8AY+Y7F+p2/1V3dJLoRdYJxu1IyuSDtwme8b6BfjJnxS4WePp565Ss+XhQ
cllGKN51mQp5tgAXPwv+575QdU4CVekFzGNP8/YEbb2ybjrgrHRxgbbMDx7Akgnx1oWVaXifusTR
RXgEZ7Llj4ttEP/1KxFCtK5OMzLEJbyWyQY39v1dvI+2CTn4NsoaUvWijCGipBBswVRBzxQcPlFL
uqW3znz12PjnXuOjtplqo6+Y5sjWgPzPAFUWTizdDInjXbROrQ5tJOD99wpZq8APEqZ6eN0w5VBb
Fghp93AqlPbF27CzVz5dGI1p+S5cgrf5LUW4ci5r27FnoZG6mep/jPuy/91wrWAIBM/Z4bcZYLBO
8etKzYXwB6WTXDVizWo229GbhkmAgi+mdLLOcBcQ3lKezQOZqyA2g6scCGuYo05JZftAeGt9f7OX
q3pqClBpL2oytP3hCLnLf5SLUVzpjV0aLv6POCT4bckvYvI6Ww4YasbUM7a+IqIfofBBJqlSw+1G
pTCC9tILg8mP1L4L6c9Bx8yQ18iKd1Xn/dS++Fs5ViOgM/XALrHdQjmCusg7ymNSgVMEma4WmVuo
rJXUw29RvSCWIMGDjOrRVRG8JglpK5A2udETqhGOFSgdjdqlz9JASoAg0B4nMe6waOYW8Up7Hxap
5pVU59Dy6fRu86VSasw1ELIyeuVfDvRmJ3vHV80/x015Rg5WYzlH06iVrow9TV8JGCfg9enycP/3
CbR7nei9Mzm2T/nMdTSYWdgSdFdSPFhvSyaAKWhFaDAasNR3TXhpB2haIfNMIlUHacYxbjR3M3Hx
FKl093hGJyY34jqnhPHdbmdGfbfH47NluBmrWZI9N7Vi1SnwzCZ6GzCEs/zZO+uuca4HQOgzoLdY
1mw3zHTtgE22h9K0XJED55NptJIk3ytBz1WKhS87oF47tOcNSNEe/31oFYShhzN8FJpTebs0YnL4
6gZz2NyFW8ulIpgelSlbUpKH/H9mBNw0KDaAWuuIw4BXbqNkIksPhm9WwljhYtV+Kk35Rc5bba3d
VEsT616PDx5kcjUz1YMhQJpOuAwy+WXf//Ox+vaYDWgPywD9w4ubD9Z0wzjEy0QkE0bHF/KitCV3
AHhkdfit6xM8xbD35Ze4nSgEBrMW9zgzVwnhAQWEcHtDFJBbPsAFW6gqHE1VKHSQfTmlKoJhXVaA
aVjw+xBifoMa4dYyuowzQrGqMjural1ZeJAJ5wDnHCD1tjzDrvNkCA6VBh7lOKQkXOaFSG+XYxI9
mConXLWAnEJcDJRCdityc8V4rl6BjvLXFrVVWogII8Ei/Bzr4misQK/O9Mh0d7/O6nVfIAwG2Svp
7km45YZhiYJxmW6SoeN0n5lAtlwc5bfwUdiQSe43E+ixuv0Gg+zBYBzopZgR0FakxT8PnslJoGZZ
02u+mtTG6aPMQGKZEdrDpBs3TkBYw5yrIgSUSdmy4szLPgVDMBjeETtN/rTF+QzJxVEcQ1sYqhCS
EvO7pfXDS6FxJjbTm62FfoJ7g7IFKoCkAlP852w8Ym56UQ5DunkGAdv4PJJZiB3YT72gjhf+Lhb1
aY3srAmWSSPr6yxNv+y+9Dj36Ovjz++0PFTcnB45Tgmy+OflsTEC+He04r7nj9RAVmo2NewyJ35n
Q+d/PPu4QB1g4Rsx7ArNgMcy9ezKDm9qAm0ffwE9v7x1BrcuZOtTrb2F0r8MiEwJhMzkPuzNZq45
f6fMoSsIZTMr9l3jiPNFHix6juBqHiOsFPorCvNU4HdxkR6Q0ZV/0fnbr3TmYPYj15m3D66OyDFi
1GTqZt6x8+OOb1EtG7IxzstclJVJ1WkHYoV8Sv6pHpeT/i9RwumtTJTJ4Djozo1dpHRdAEmsH2C4
KypoVEKSgw/dlH0JGRWDJaurGDt/ZZP/rOOk2G5g9n1ntuhnKgwen2rMLfi1QywVG9mq5p/BDo1w
RwR2s1iHHy1RjS19wj5ttgjIzG6De3+dJh/dVDIOwYW/L0NT0F/N4iBQTZOmpbU0g/kxRhr0bCvD
SiyqjuYmfptGqfQbeh0NHceg25JJI3/MecstwA+YxPpAfkTTv0fzB8hbh4kyeRRJbASPjdKVSd4J
8BIfDjfrfyKq1OLf5SQqfLL+BAFKgbm8TelAqJqXllmiov7A4eGlqh3Zbr6bDKIm1CKk02B0Q+Gy
baYoFeuZr6Lslla9uwntIVlI9OYQj+442jnLF6kh0/128/Xll3ZE9dFesPdeXWev27o8DvKRsvJ5
IjfLqvKZJvkZLfh9ngjFKio4bOPoikyMFRnGJFpbN4pQoUmXVXAfpI9WUU66DcTMVlWhJ/GEPltN
wlFgrD757gqqQaXJtnwcDLm9Ye+uDeqDyXPqthWPKCHaADQ3EgnNpojJFWoyTAulj4BVSoKn5lRs
WPmAotcz/UDB4mhO2F2Zhli8/PMlYBHY1INcrTMo4cwmm48jzYWEAA6H9K1xNu9KfoDDqkrclg+2
t4yjaexy65t7DG7080paz+icOGre4W87p2tXrlI5kXA9P5BQNk4Fd4yCwtnq3fh0x6dLopR0Bu1C
olrORo35YYjejcXk1w+2jQHTiuA8GTsZSd8kVOgPHufCZf/9CydYWHwDeH8qVw30zH3JORhKaL4F
+Ok+2fM/CaKxxT1S9D8zLJAA4Sw45owno/UKj8T5JBJiIU+6K5fwxXZyVROCEF2husP5Ip7Tv6I5
XY6QD5yjnvF7A3WHkZ/kBocJNBa4M/uGS0FawHNRt7mCaNyo76XsH3lBeXJJlRsSKxiq1yDeqpoP
3Bi3j4QYsfx26kJqB+DPLgNPaQEC8hA50fumPjvJvClVLABMVRwTScp2rT5g9b0cIZrm86OwyJkZ
TJLQQ6zDVwI7fzpkC6eD76I9lEOQHZoG8qA15T0S9wuYWFkQFzT+49wY+cJpyaehkK4jLtwTk3cc
2LhnbGcR+F91rAHDv7no9d1HhEVV/MuLExVTx6YkOvUKR6DyLVjRqCJdFy+mOqsbfHRLE7IMasTK
husHEDKJXymOGWmnyM5f3QdC6tb3FCaI584fZT5N6Iw7bJGJyOpt9V4qCMkmBG+hpSEtoAoZASoy
ureW0ST+CtxojVj/0jh4xDxDUGU7juE53O42ZjaVi1j5utInsGJocIzWw84+5QAYR0tdDQccBOHk
qMqyzaSKuSmqlVf6RlWads/xWDdYxV3JDZKdtfnOcHTTOpGUiE2lj7TxQ6Q20ILHdvOC9g5W+Vm3
SPFtQ7sQvsFIZPrAdthXalT8M4YwJp9T9lRbnsYNoLI50B/GURxDVaMguwU0JOaovsDcabcxzAvJ
v9dJos9NzBpTe/zi260H4NmLH4/V2mag5NOGYFyFQgsnc2Vc1OjFodxpB6d1JwcKG6+U2c94hDkk
OxknckG/ZAApaEXMKSyU2ub1vrpNUWRoRQt44t9hN+aJH09RpPgztS9oGA/4WXIZ3uSe7DOGbit6
HBbDg1NKaLsXX8CdSBHZ8FiKZH9O3Rx4aZLebe0ysHLGEGgjHWT3y+dX40eBqz1Nvpsruy7+nZrS
y446gI3hW/Euc2jMqXZCvz0sHbY9tlEtpnYZX+kGGJgussusNg6ocxZxhedi4HCDHAhTaPVwQLb6
CATqlWxO8wMz4g0sSleUDmBjhKvc6Wqs1ObJ1mogySxEgDZkRJe+LXDdi3VF6XyZpWbAndcdQs5r
N3uuch5oJVFOORG9eyqVvDW0TFDKGIaIw5Je/qevEWFMSlLoaiGtQ3yAjBYu5f1f8FQ0Ae+aj3td
3Rs0FvYm3+3wLj1aJqHGFxkmKhi2SlM2SgwSr41Cs3bGHxqcaXw6zE653YSQMFbqgqpehQCnhrY9
WoBBYzngQl5t/5Kgjw8pyyBqQJ8kTB1jY25Yhsd7PseOhjY/epIU0F/ASCBgqOYm2bKFIwrbgrXT
ajzcgi+puyXedImD3Eyuyjz0kSI+6Hdo5q2sfJXZB//YOhv5dJg3jJJr8HQKyig+IcmtVknhoazF
Fcni2I5GWAmPPUgATay7vwG87lU/ZlWI/LR9PvNtQv0Bqkvxpk9o0XTVh1bC5mbKOMTKRUu21/Ic
RB0ZItikl2yEI1qQJg/wsLWDd8xFUBEqwc6AXmQaoERYlpQQoh1VBc4uMdSAFNLiqguvMsKs1Gzg
Ktf1p9EuRA7rm7HCiUwDI2/jjXk60dgYXW/wHAA8bhHOjdr4GDogpsh2ZmusQgwlhb1rC6Mw+iVg
VGXcAPxAr3oSHvAzwfcI3TDbxd7auYsg2ZbyxadF5H+/5Az8Bm4cylBYIAF2bVZcHH4rUTQZzYyw
NpQzRv4d9UoKTlSVuKaO7HgAj9JJqMib9mH7nJmxkCNW7bEezt6TC5BgcKSKEFluFd8YS0ozJa3d
kgISeCCq7d6A0N/bFkyLM7oojydhdWu/TiMyww1vs6bZUPgmCWWjyVyv0jTAgnbdPDulUSbPe4wO
i4JqjbhB8zJf/h4McnKGLkMmz4vTNdUv6LLKqWyPVLHhKi5b4L+nGOpoKBTkrbzDFa4jlO2zwHVa
FAvEIkaJNLx2sbQRIASeAcsJaTnVs4Ec6GldRwdL801OoJb7kDb1hSMK8JcXz9uzLIwtTGnRkGzN
tUL/JixkLaqGA8SjUSnkVUWMn3x6tRxAYpVx9fAeddsgTBUwQGVY0kEnFttE5JDW3DFAGdSRENax
s6pnRJ59pgNA5CuqPL7PhGb77/9bwqqwjbDxEC9eB5R03BI7SVp2JtCZFxcMwKrvaQVhkhJcolZh
xsjA8zDMGuyE3fuzbo894d2qzm7Yy5L5FERPXqFjqR8mBCMPLtxmezPaZLszY3QnSpOwV1ywijVb
G6mn0cGOWlI8HFoZKhbMIC2zKy6E7LDdniZeVR5uRwXPzqzORylAu5p6nh+MNktj0p7q+M7lyIuK
NDGbnOHxKAxzpz9RxoxRH2eT1NJZ0D+ZX0cdQmoox3oQ5T8RF1WnQLMhFpgfFwXtL6ZqYUeAEt/Y
zx7ir+cIG3lopgwW5JPiqFBwYhGqZbH7LkkteCc+yKod8W0M6LKTdKtzGNe+aUA3JvU8/Paeox7S
u5R5BGwPD+0RQPS5rGnj5aqkbiS2YBNuEACWb+liALLtwpgmCCIbdnL0o7E5pL/F35mmdTXiB4GW
riCZ71G3sZ18jaDcbLTXxAVpVDxIdUjGm23vQlvTqedz4hb1x9TBkbSDhnA1PAPqbCu0Js3O0Ka2
e+NZxU8mWuG2DDTx8vS9K8sBCZSbpCRDRpy+il+bjwavBqf1dn1t3R/dDiQd9CYCu10SzdIG1xmy
mHAAETfXMyDGMMl2WL5wg8CaCsnFZZwFujQjGUrJbxzJRKvuarEMx/g3wYqs6Q8mqbP0Emrcsuej
0wko9+mdbnQjrT0vW8FPDskTNyzl0PQTvb5Mh5Ip5nPHCSGhnorRXG6KhuKOlvwFLP+bbNh3G88L
h5NsqFJhmQzQayxDThfu/YI1YmHPKJDAyUKYW/Xs006RAcrSmr0DjfmyED8XRfo3cDZtBIB91/2w
o2WUNYvy16TyKftjE1SD7JG4wSS9dDRH9OjSR+Cf2GlR1DqFPRBhEcvCZgB2miejCJect93Ao+uO
OQ8yPR/JLqGDj/C7uPB4RxYhEeTlYE8VLTXOs+0BEfK3GIRPgqGaXvsNMf9Z/sF9vbjA27tUXIsb
jeLRFQ4W1ISnQ4dsbmXkJtsYE7INq3vPw/Z7ysF0FJC64jplbZKPS0HMjWQppzFLolHv/pZNR+4W
Kpn6bRos/miMXQGAs0Q1R/Clu8Jk2j5RWKv/wsYXFXEM+2wR4jN43u/KcPjS5+x68CEZZvmZcfZB
4z0dSCASOFgC8KumI9Jtgr0fBteAnebRfyAEvS3NNc2CCyLszdA7B20elI/qMX/wvcw+i+aLkg0D
4STGF3a2xnAq17Q6jSeljeSZuG+C4XtJJw/w83D3fGoXnwcBuYfH3z1INKYhmxbyOriWQAJMgG77
ZrFUPSK8E2UdaxCaJjyNLPoCwQOm3Dhjhw4yjqX7wS1NACUYdj4PH/FOq1LM2kITObCjH5v513Mp
GrfMHyBJJEWsVB8BMWVvAtsAzOI4PyFykf5nQiahuTrXfRSBLsdirCqQ4wmWBmiC8+0VeTLp3Ogb
vKlFrCR7t3FNxyBzVy8xPjVmTpnMjf6GMs0N6DbVNYs4D88jbU+zBZyHg3Jx2D8OTbet9LE2l0Mk
EXDnsVVFnTeO9gNRcp42P5HWUGJtMkVgN84Kj0LHh66z0Lq+U3GM5nBepj/lnST2dnJwxe0ikBqB
4CNb7VanvXNCfR2Qe9sKyDUVyPURz+UOD+wr2DzO68L55vztP4WLCsaBmfiGpVXf9h/C6ET+K92W
xME8trv2L3Q/CvA92Rdpz9kWnr/Fjfhgu+j+q/KoT24yc8GieyBhp3hqfrNw4z0+iQ7ub+TQ5PNy
R85udwcYLD50IjYL37TcdglBeXyqYhyNf+fkXTlWYdePR4m3aYxZLp6QfkFyI4q8dRMV6au2qcTp
kRXAAkr8Y2fD2IDdaAXtrFT9Zda53UcdBIh/GxsddI1+p/HsYyqwxMt3GyHCoNRUV7H69gpTSBpx
+5DluR5gV93vrgeRyz29KknoCl0o1nuKtaTF1cIhVpMvrSEccHQCcIqPsNG10aXgPyXiK9hN6DzN
sX+VZIc42JpVnY7OUkj6Z48At+fxeEykZDMYr7vFisXGGHSydUonjS0bUKXwXKa6l6ECouYdHFqn
Oq5zRItjlTeTpOWcrUxNQjN3lZh9A22VuXQD4X3AQtL6YTIJZIW2GdhNMnXLFdUE/u0cJ27n0/oP
jrnSFfqItOrKxdtESzCLs9EGk/q8G5JZueQzYTQgZVjJRmX6ExlcQD40am3tSnFDzgYlX5jz6byq
trGh47sN3tiI2pEwaZqyxo8J0ieBvuP9XC8hLinoRLiqGtdTyh+LExgTnMUrT++CDUv4CpiynOAQ
RuI6r32CERS6T8TNzxTTwhDiSDc6fketzGUFoAdAMt5KSW3Mc0HhAB2YdaiI6pi7EvWcoeLwVSBX
E7GkSuBEwHk+X4DpKkzur6RaxdbYTh661ALKK+hl+SXJBweKtLC4XPLK1/xEaKwakh6Cd+87Gzf0
+FHBrh1QtAkklZXQg0yy0pGLBr4I9bSihBEt/N1CBmfPvdHEXRL1vDYag4xmKBN6MQBNdAwl+9KR
tb08zDOh7ha+BAvGyruTn/8DHHGZFqbUBbD/hnz3wvtQWMd9o+sScO+Io3n1Xm84rwKUjcGDYjhT
p1tO/A2yQXiDItr5ZmKHHuezLcvfwMUtnJdCNW6a7b8jb0FQNpJzUf7yhlCNxHnbZ73f0fzh5clP
Z3ykfyRvF627qmbT8oRGkMI/R3fv8hMa2oEny9NKkM+o08MLreqDWkf3k3bc0uFuXfL1eOHCi71u
+k3qvNqMTjV7BptRQxWb4LhmMj4e3KRjfHCvmE3j15sjj3gxMK9BWWx55ol0kVX1nSKhh6ZjujyD
w/g6BI0n7qip1I9TbGKLgrFRlmUE5uREjw3vY9u5sK+fH318Jf3vn1muro1B/yjI0imffMObayvv
xWtIqANbZQDBVjiL99dbQ2Iz7BTNJpYftfgSt8k5BaaxdMFjw0doH/zXzeNGhZK5aGGrLlUYjF+I
0NvCHyjwshljXlc/JpKMkS4Fqku8/AJfiyc1b7u7U+SymAba8ZoC4RkRH/iWug+ojfL+6B2Cs6W2
iHNCvUd9vkEedN5lrkunWb5CveDr/RzJWqKsw5dPFAfnNHW8JP3+tKRsgCUkt83ruXwBQhcCOlzU
X0krXiWKSHFtgpsJwqHZEU4GIIGYx2V2AhRTPidKvIU78cnZBvWZN+ZGb8LSh37L3H/EofouQ1YA
swXkSysDVsURz3BREHXVTGgGGDdf99L8UWfX0Q00VtjWmpOOs7eAkM0aOPisRSEbIKg6bpEWOlxd
kjmqchDJQtZCvMjrOXTZXtSLiGpIRSQJtS7JlE9WKL/wwlY2D9uZFqJTynYrUmU2c8rVYpNW5Knp
qQ+4P82HwMWzz0LrGxxzbIXAz/httJprab6PrakhxaKKQAsBtKMXFNPjExRPK9l6UIhs/wNzgpMs
L8WEbVunzR3ZPY3l3kdQxxlOdNFhMB3LJkNodTNDhLAYW/BUzgTvXZ+gZVln5xkUPksXWCuxoqZM
2c69knax1iMxsd80XmVP5GH/pp1nyr4NjGHSb7JzhlHhbbZ6/RccCBeR+9SE0mffavz9eVNE852i
8QO/QqbPI0TxH5bEA82kOufVLecXrgrKBlYzn/gUT1fWvq9Sfm0tUFcuhnMYnVbr3oDBcCd0cOoZ
rC5fdUdOXo2ShE9uoCNk+Ciwc/g3UQckZbxjNHbrRp19qrKPLWqrrDpkpc1UNhhEQuAOfQ+P7q45
QIhWuEv4YlOGdEPpt8aPiQvX2JHO+CUiwZrHf/sghJaSGTRMfAvswjPlrf/uuXew0IdATQ7kltGn
Zru4WmdZHncAjKH2HwfE6c1l+mbEi8Lqnfey+ANMJTc56rsqq5RJ0CtH7lSOLW30nYxceOyxAZEZ
29behkyzY4+vzuUhiJsPdx4jV8uQpJWX5X1iRUseNE2eSS6miXIVzdhZdtvZyTL8KSdWII070nTR
nb0J7d98rq4ZcQ/K9VnxppFNgcQacev3x9U12Wyfk5o7qtW0eaaPc3RVCFQt44ULD9NEI366IYm8
xqCUpJVBeum5J04QyyfW9vKQyuAqU5KV8CadZRvvPTfsdhS+7aB1dPfvzIfQN5/dUz5k7S5tLT8m
eTb80TW8aqfcwxRYlceDTLRGXJF+TzHV8comuzMEhwSH5CWuv5ATZ3m1lQ7C0lg3AU4ZKxn8ZDU6
DST4llSIbE6RX9/fJ7hxepXho16sh4vhMiAESPZ80ibYg94spioSI03dhOxQfEHKVWoWp1/ZcfLW
BcMPJe0hrYdNxEzeMdYhb1NirV4uIy/moyeTGoIgNpGEb+2poKis3F5u8kuw1k29H/ar66Ce3P8J
pprfMJdE81xlNKw0PypOB38SiD4gu+WSmjxtXYdCNzDD9MyPOYG212AE+WatjcoUmSqWW/B6SPbC
i/Pg44bqRnCvJ7llXR94PynHcJ1XDP40pZpFWyb/jUreRYbempCYAH6zfsVps9HYAW1+ESoQfYys
FkaQjo0BIEDWoZpgwQ27eC2IKGn2vugsZKXSnkQWpEtDPN4MvbFoZwOPu/bavsq6PtoTuLfBCheC
4XgIwVDXnhSXQ1ViaRVAmN5b8MDz5yhYtdK0cGWLZs2B4syTKt5xy2n0gH8hp6F5/25mKLrNIeYc
K1KlZNolE7cSI69G1Axdm3RzqnUKLvjA98S4P8+7sPmG108biHI6lL6Xln5v9vSc2zowMO1bgpgC
WUs6kewftaHWS6Z0jkSDk/+8og2OSea7hQpAs5oCxoj9QjIUGw46xzw2K0/Njo74p5ngrhUe4e0o
D6Q8oNDFYL8T0CcHLzy4/mJiOD+JDrUH3CxDcBK/VqGY5XnWqVNaACH7ezNzOQU4VVBiXGH0j0ua
VpoafTus29vfK/1oIafSnrTKdll7mJVzg0J7ygV4QHAogiFkljysC7KtoBnLXCWICMmCI+eJfsWO
49AFuLxUcXpGIfTMbvEASsMsAtvmRoOAc5BDBF/qj2eErabOJDlw1aDQnd0yOAezrIOdoi3qT2mv
rxEAWzJRCYPMTuVqkOZgTM/s3LwfFoDiqwrqb3W72SE4Jy6OQ/PSbtJu3WFKWAIdzxCspmM41lUF
XWkfNeALJC4JSQmTwPmeRo7goNhqt12hmMhMJz8hLv/SxWuquYno69uIvJkDPbik3jZFOEVVYn2H
nMcVOiulDgEbk/2hLZsMOAqADjzRM3Pcobd6NaK4Dt6W5RJGBbZ4D1M/FEEkl1fA4Z6VMr2cfGw4
xaE7V/GctOK/uoWKSFseDjEfA18RfD1quWbdHsyvK+tWX4OL2YfSeU9TbOiaJ22EZ5He6vzsZlMW
tQ86Fj0JURdOrZqWS6SeGEcrt2dUH85cy/V88pSZegnWGtYXFH8gfVpEnANq9bgCdg3N/WR4Ih8D
BfRDbd+AhQCbTVHtpJPMMVMkoBCOfDsWx1SYlpGGAZ413KYO7uPKIHWKVDCk9V9lbcsecY863L8k
xuq+vgn5QOcbXVIyL36cBCwhUA81L/Zj4XA8XENbSsD4hZJMJlaMIKVbpx2wJPMwwNdJ27mlRTfI
jvLuaFIW0XOkiT+VaFeA54VXc3WMhdjPV1NA3DyhEgaUBiIIhhjD4iWGsAweWinWNX0EoHSwFzPZ
waU0TVyy/yTRO9T+u5/lP6O3pjMolGT673LZJSU82Qr42vOZTfIsLMj6+BEYXbkwOcZ641/Rxv8R
vscDDn4yukBEIKB+jK8PFi7Ep+TJHI/XQqo4dtqANQ2E4tFUYAsNFrX517scc7FSOnrs+tqOLLWy
rrV05I9Gge/igjPi/dB5P54XcvWNCPiUjo9sj8bsKVjjp7P2949/YCl/SncEjJUILkh/uXVoND3+
44o6y2jCuNoEY8UZ/ESoP4TMu1zg96G7OF1CeMqdQ2+pMZulvDQWojLPqoAjI7XzIf9lyaikZoD4
3t4UmnKhpGrvWayRoRXWCm8BT0MJl13GHxGeosIXPvCcx9kjMBixYBs0Cx1osNYbkSik2gWXBenC
ZxLSfW469r+PJIdWQBae+kZgG2L3lQMMnuxtHPX7hktT3W57zMeUWnmFZY7yHWYGKizqbTfm3k8Y
jRI6F0Uy/5EXyHpRVTwqGrkv+E8qbUIkGZm/trtG0L12Nq5DHIVmInr5kz1tUZDXpbpskIlm1wi3
A6fpxRV17GKCU2ydMZow8n/4bDSZYSEx9oCMEyL0IoLNzZadkEK01PJfLwvmg1+9p7GmI3viEu8s
db9rC86tqDf86OACFdY4+VCe75CHQ5g38JGmDm3T1TqK60dcJZj0OwSn2KiO/fPQY1bJ6J647qIB
HSzw+gF5NErN1MZXf+IXunaBhg2Yopu/rbBOasxxdY+YdlP64cZ7C4L555TjqQwZd5eU0w1y5cMI
Z4hgZko5fv107B8YMgi2e4aehVe+/hIi0ruHBR8vCmWNkJ5GdMIX+Z3CYuH6oXS0gP7fO9G7Q4IL
XMt/sabX0qgcECcV+sneN4eXqpVr3onby6/F6kvg545jVYilRrdnw9ndJLHk8/3VsocJl3BLNx9N
aR6Yom07hZvcY8CBJFRoRjVE4GTRudcnC7/t9/rMx0B2JAYQv4svuMpK8u39tSXrkTienWagoAxn
3OErKnt9TP1p6sKAJdYBWAMSCAQPtqLaqaK5ZOBsHkorvfmozmmSxDRAOL5Y5FrbZb+50YbwQz62
vX/pIC8BM49nNv6w8yM2tyVw8swDgQsUJ7VLLkSmgRQN1KWjS4nqGoiHn0glvIZRX+5QN85FNERX
qnT5Hv+p21AFALEOyBYFt1g8oLaBG04rgwu5QEE4hQj1pByk1KpUIXDwv0NVUu9tK51OlrS7EzaI
Nzw+bAAD+quuQhPHJSnle4k3+V2WJ/DhcVKxm/dUy3nkr/6GAgUh4tmIQQpYNKELPrAZOKfeYHH5
dbv40cQcUlMfZ5AMKQDkZUMy2dYosR4ZXYsnUZMV8UJ+HqnFdNSqZkXBV8Bvue2AXEXfaO0Fnj9n
NT4yfpeUCJXAfY+B0DnYKctnI8CJ70oEmmzChjHN57G1bJit5vYxIkt2LOXnRiw1djkPBuVxyDDR
Jm1ijoTzU1GFHO8C7GRA/R3hQxiOOpCdFWzIVZARcQ3iA55f2b+8s8OlBxQ8a9lEgDIdMJUkmNEu
tdKuuiorvxec6LtonrxJ87zQ9z/JkbBLK0/m2hKt5CZnCMHLSHEYi1dAsiP1bY81F1uioTKHv+kY
DPv77pE8HShjIwPd8rSZkrx3Qwv6D0DMUezR3p+GI7Gu/4T1aX9h19y93wR/uBa4o02TyJcFI7bf
V01oiifj6UC1LhtO/Lb4pyxFs9Zm/Ke1R+5LZDHP72wWJR0qR1rEljjN4/fIC8afNCJONxkUvj2L
ETVK0qXHlbJFb3seAUSZAWuswWG4QgUBazlXKL+o+CU9RpMai9kevEvXeOSMR25HfHmMvUrKJ7/1
wVk5IUaPLWlmpvGRcAa0GmqVdIIoUFr58gvQMhkRYZxTwFVI9YaxGNngZ2jC4uaXd2F5sXFy5SlB
LO8E2YG0NFyLfz5V4Eh2gO/5HKduqvaoRIljp0Tcgf5HiAdrNtme5MqM7RUHvJ/AYdUGovL680By
6L4iSSwDnZ+jjGIMm+ODrzTLEP1ooE/ACgC/Emaj3in9X8md60mCqpjGak7ClnvGAuN5CdWRfRNO
V68ak6fFH47XQ3k4Np1kghknfHKhOeXhS4hRioprP2ONnPPS6aYCSD7Xa6sJo7eE2rZIiu0UZgKR
UtIJtCpI+r2y/aOu9+jZtj+QiMoLeo1x+7NYNyZ3cjQPV/eeYHYOf6S0iYYCS0iwr2JUvBOz7f15
ggFjeIZF7xRxZwMrn+a9yIq+0/NeAIa+uPldHqq/Pt36JTafPm19bpj1QI64x4B//I6uI/vur0Tz
myHh7wcnwgv5YXlCyoq46aCD+wgUoL7G4REUZnh2E9IUTTfpxL6XyZPeU4kUkVGaQyV2QEVfPFsm
miauR/pAS1LgIvUqBgtavUd1ykw4z2yNgQnPOqd3hSnZ/d87RY3EWOj4WepbkGSa+ftL5EKLsOj7
qaWcHEHxOMm0W98KCI6B98CzbGlbYAX+Xcnbv1xkN3bU6ft95VUgJrVFXGpAVDs3kWFvllaDvpCH
oRYqmFmXXu3fKyFH3bzCSo4JD6wU5mvWVvyoIKwp0Ksr3fbMX5J4PKqPswCduL8FBb7wLWAYKmDX
uCgdftvUh8Ekwn27DbmVQhR1qyUvloEpOmCDop3FSGBeOwElXZ1Y2R0F8YK/KIh08NO22FQGH6TA
BM9KoqygLJEjyRQcBOes5/+n0SyvZ4cADMH0o5tEeOucHGXjlzJq5ql+8mIzUAfz/UrMZ2xOs/gF
kfNAjY1sdo7LiPcF0SkyTRXxhjayL1xTOVHqeQaLPOu8/E9nR3T797ugDK2nnD1bRU24w14LRTCA
pn/TlM78LhtntLzkbsjOtaBNsxwtptRUaHZ/rZGJRD0k7yL+3LwTzuYDHNWbPEwkjSnyocSMI9ob
dtmx2+uBImQ7nrt5U9bHuIXatXeAlFcbvzfLpuALFpaRUSLhd8PBcic2RJjicpl8pj5UN+FIohpH
HRIe7L/2l1z7t+0QkMSm2HvuI0hOrvT41Db6N4hWbikin8J52ybcPQQe7sVhRPyxcslT56cVDKRE
Lb6OvyXZs2zSd44qCUzG7BRjBLbG+fl1t8pJkCXDCk9dY05yNK9ytcLlRLIMx7hLm0fCNvwHkax7
AYsTT7yipJFfdSBEJ62P0nQn+oi0A5WuFDczEKnEKY2K5N3bIUvaypIA4BMDsYNmG997JLNig7a0
IlmdaH5vqzOy3NelLH6IhO+XY3n1l5lPO+M6stXy3jlvFf9q9dPNKG+1THjrythDZieR79SY4Wkm
h8jJNhTQL/YNNUrHWhhJY+ClLhYgzvFZMvPXKw3f/FzJJcqx2FQusH/osXgmslU0AegF7F/O1aDk
5lzF2CcuQbZu5ZZ9LY5dP/e5/9CpUwjNWg69l2aYeWsLcskGroWWeRGti8z7ZtCCSbdpiARTeoYe
3KTzu3wVr9aTvnOWwSz7Nt4xVbrwzvt32ZT7xRMzlhZQGZmll7kq6ekthMjOAqz/1ITFLZpH+SNC
VvtqXE52mf7+eIIApCOj6W4RlgnuY25YMgt4Iz+8yhP3I0oqOlG2/hK6nWUbwzI/7bv5qctWkvVe
Yg3nrmM7MSU7F63zgvJQPXfHIgW4f3m9T8g43cpSfqcR8R+NatQdXe8u2KYsw6ZOVxSCm+Qg6yxc
Nh14/YOMxykI7UZg+Iu0corQhl5ACLNS6Kxoi0biKNlq6GanSLbqfaIJs9xVSC7XOSluyRFF7rHO
NRNw/3a+7ImxvKqS4kK8+U7mH+gzhRez36lMCntne0Xyl3qg++bqI86clpi6rq2Rt8T5ianp/+Go
k8REwwq+tT6Ewv63ewJC5GmcKN1R2scPIlYLUay7v7Y5+GrqZ5k/HrMzbUuPJXlMnZ7hU+PnG7vX
Gufc3u9fBkbCxnCy0Gfo4fx98QDuOMcusP139slf4ckmIAYj/vx9f+iuGt0McRbPQmKS+FqDxtMd
gLpNIrS7Nf5hFuIHD3llU51aj5xIubqZgC/m3Ar8wlPX5Ge4dUYsENed14+RmrFHqEjUd3QihmQZ
+ft7oU5Baf+fCB4J6TT4YEPQ08MMX1MfH1pYeLw9WdCtIsvLf7K0Ci+wEFcD57YgTRR6ICTjy8pD
zBNU8HPMDl+SgNPOy65nNVYeaFpsfKlP4XNujJrRT73WhVVQxBaMIzcqmMJVvHurYBjvKNAMqEXl
+2Lq0hOIAV/jYtsNS9989cG3CkFe2ANLiGcR8NEIcIyGXzZljTylUUuLeE5vBvdJsqrsjW2LurKe
PDRrb8NRU1ZgnmHodpjki9QKSFFTgHlTDM5kzDxu1pNXI2K9GEYyLV1QG0D5DSFOV3IAsbUZs4Lb
0HDxMkVzN7VRTgXTAf8jUa84ymQcQhU7uFccw1VKDKoRs2h3UPi6ETcTZY487W/Ogj4G7pE6j0Tf
PonbT/3zVjbmi6atbI07/jZE8KensXKswpqWPc16Pl2oCUKDW16xZlh75PB0yk9mhY6KgHWcwxt7
Bm1JQWdX6rhpE789YBA1N7f7/2/uipzf/9JbuvzptqPqsjE/HDBVQaU0gD3sJvBPeJgJsGs2RAK7
T35r7P0bZ/X03Tudx0TvzOSsv3BjRXrUSjLJ5Nj3Q9s4KI89S01DgikkaYAxCXHZqRkExhbTkx2R
ozseMGDimzxLD9owPMMYtZZvCA0jIgZ4ZaQn15wp/QfzbWA3TjKCYzmGpbFY4HOEGMY8xurKrBNQ
/IwWMnQ81ysfjHS12oZQybvKVWbudo6tIMhOGjFftU22ux0xk5fMMm4LWeX1FI6iP9KnM2h/egR8
yw/Eh37kGe8YbbQp45rPy7/2znSi0awGFXTQx7QogUlLfXKdq0aqzlAeNHBWDX6UcxFkUFd80pkc
N4MKUZx2XfI1jbVXgOA02szXn5N6b+LREJCjsdBxeHV3MeLbMBlb1TAKQdBT5PgeoLrvvfDhvZv6
C+G0iOKZUT58qGtwaeQlb7XRYVqz7fQqBKRWlael6d4/4IGTbgruznqeVUyqlA7WLrZWn76oOBzT
t1BdrLSi+pZBQk+3dtvl5Y53EUNKOIRUpOr+NyHomZrER47vnDN0W3+j9OY/rRF84Oo8zVKIZksL
GC/EDp+fMZawy/kxc6QXI0jnmlRiSFsXVHV36rTGjYsQ6kXfqUeXESZtB1GnbcdPA1Ju85jplKAS
4saByJuSAOl2xhS0ckwDSxm/w+uj9nUIkF3IozRtwQakFY5ZzwNEfbpLKYGeiiYkbDmdS6dpzqrZ
xhqYIH9S4J+CSEark1U3Od5TqQrMrFTOLqiHZWpPAaamZD/h+aakeisVq+DM4CbiRp1oYsxe0/yU
ygNmV7tYLd0bmg/RXTJjivgYXZxE9Op9DHFBDXx09POrwkWa3MwJfgQaP+UDW1NkPIgjt4bahmx9
6SmCs5mlbRCPMfB1+lX0Ym5s7k302c16lcciPGvJHN0wzwSvgF1oRgfsSUWr5ETTsDXRPe9QIkTk
Fv8tJGspINQa6IUFAHhq9IUVrLo3+nY+kyCmioEWieVfl8tylSFpi4a7S6/WqBX1TkDWNbzJOu7/
ybcT+p/A+22cl22KDPRfK+SOaijxXodq/W7humCmIVRLkuixsfnfmHD7tZ7+Vi4PYq0U5WFJTf2K
Q5y49yUD1AvB3xnpjFwYrktdHNXQ4nKPw73cKmB3AvNSUKcENPj7jPjM/sV5kRDAHIocfvyEg+vS
bPSOu7xBwXCLE9B5Kha2zQQ2dyVuuIiDtkzVLgTPy2RCOx9gIApwT2lIV7HQ+gxzpwwcC6ybXGCb
LpajcHUeNZBatH/xWZZNxnyF3tvr63ltiz+WhC+PzO5k+MzV/RZzyRiKv1Hdp3g97mX6KXp2Soj4
hH8tH1rSAf2ZEVYpK7ahUhkOiqPqp4nCNnsOIyUskG3nIk8F5yG0SmbzPmXE4restO+yQEDWmg8h
DeFbDXySQRRr8Y3suM/BbweOVUdQvQQwy9bPXKC/KI3wZBbskTEN87V7zf5fXvWLSjxYja10VT6O
4UcBuYjFRpcdIZxFm068NEZjev7N9LGBIqYPGvdClj2Om4J9hnOGpMaXoE9ncAQ2bkK7OxtuYdLe
A1Mb5LTCnw4SjMlaAj1iEuuardrXGupFmM9wvwWyXqkYR8bv/7eGHf7l0jXl2zMqQODwQsV+YcSK
oNThLcx83Fsz/qFjt+AOB3z1n6Bp5ZXmcSC+HPwCSC2stShlbgom5NmuLC4Wkek7xgb5f5kLMWb+
x0tY8nF1gZMIgeGkxbtHXarrzTqcS6no74WMfsL2MMFAYR5jmayHKsbJBQ1P4dXKPDj6097jxzmC
PP3iPN1jG1fb9gvcECXPFHkS8WFCQiZmv3xrB8SyFU58w5HTAtdHmloo81/rKh3DdK09YRFJqqgx
RWET8MRm8ea5Xh1kwlK2KxNWEP3CbfOoqABH+BRqaqOz+24jxiYxG+ywl+ysbiJYZS6ktC0Ea5bF
GCQFzizSAQq7i3/QzeGmt86+hJmy9xv3/MRtqLOIyuWrcCJFLnmLM7fucOEhHHT6IUUyTi+ZxJIu
v6OcQ7HCo5vTpL8J0tnkR+wIN9yOtqufXaV/76pv+TsuUdPwOCMxorLJdebP1NZH+LjrQ3Ug6KNo
cm+aNCkxwMhGi38/yR5AJgGE5ocnRC2vjDpixZsqEB4+oclvpxFdLKK7cujrcU8XW1ORKhzdMncB
E9jk/IFB9kcrpwp41BvwfNyVp6WOI93TFii4JxWEbY9y6JPlO7Ke0GsCQOE4YPRwA0CGEfML/Fu/
fUosdZy/+wg1F3rZYCKInGDla3jmao7cH9GpXjYGGIlTzyrpJxUHcQZEOJbD3+YW9uFjL2ibbpEL
/p2kYyDuVe9enncd73x3EAhcADYS2pEc73uB46/P8H1VCXYNyGmY+G7ZQAAeU/Ryna42EPJuZ9Yb
kEIVldt+A7envmrHW5B+DX4VU/Qds53HD11Z4aphMNflGtkCuVL+PtgTJCKWSDT55vbUBvwkPe0R
03ToUKNuhf3Y/x4nrzNWh1pI4n+VLDbesNh/SRstZG4XUFGCwsey92RYBjDO+wQOP/YNuD6OdmbZ
jTWylxmnESJ04T0atipOAuaFKU8ytz9MzjDVqNYrMSyP5UNubZFhu/aMnDqEjQE6rBF6kVWRWDdP
faBEHSTxAwdy5oYoXKAKtLBNg+BHyNk55/+7/uKM41AFx+v627cnhKsG0br2uNMuGErv5MoISY2g
QNyE23LAUppcj4DALVXqICDkjFLIJJT5JuRk+3BpsV1W6qJQzt0vHmgXMeKxDGkH6eRRmHr4azS1
m9FFSRrggzsM3J/iqTEFnF23T8JGiI2EdQnUS9nziw/QyWR3/RQ3snmRrRDnOIPoV1TlIM9AN+/6
2AtgS74tzbOG1IUiCKeut8f3KhwculqHY0AT/QBMH08yINEhtVbml3lx+Zsq9fUKtbR9220YSe27
vqOcvlVNCJG3L2Puv0bxs2X/0w7N9xkFa5khoqnPY71cLE+AC/UjTsc0H0GyHdVmhtN/XtgIlImy
hRqs4reFrKgLKCYjKLANTwjGDaBoJWaVQFo89POuyqxE/ot98q/zPkCBqmo5TVWAkk2rdMLa0Tay
F9BBYVqwDVBrjtw8vlaI6Wpz4bP38VLZc/mT1VXOQhVpgZdFjK06L/O7g0fKwFr5OiExPmAXnxaA
3q5hCAN4RrDjMt7Hp2ikrWo+KjOMzQYCyCod4EiJ1CwZAXktmWwnIsdUhBR+RNjurFwjqQUrOl5S
cnNT5jbtMY6EPNCL1AeNgoCdiSvCtqGiCPmPDB2eiYN/qII+PBx9VfzpQ8v+k8HzjXKU6N8iPVLK
pehoJZ7cYiaVrWIvlcw2SzCjSbPSla9nkdfnnf/YiKGsurxocbbCAqo74pntaqj6OXuKpTnliHni
ceOcO9Qhx0bmup26qZS1v1t2ecw5qa+N/OywM0tgWZKOyu/F5fKZVYo0lX7/d6WNxLZSFhnUJo7W
LeOLrdTvB+BevxsoGM5UKXOlmhGWG8n4DoU+kH4SoweH/IjVjGbBfO9sQkIOqG9qXmRTsoKBhk2P
89+TsPupti0Yu8POjwAvn9eCRoB2t0oIjPJcBIPfviePSlPoSxkqP2PPTfNcgA1GsBrocNNTnd7V
qSq1YhDG5qu3RnoevKjgopFeOFuGNOaGqz/Z3h22TLxiXJfkBDvTJnG9dUgMyd6U0wGhEuZN+X4G
cUgLzrUWOLhRRGn2+jZv2kBe0LAKJP4W+RBAA6T+HBTm5qEk7TPjP0uKlt2tSlj9oCIAAoUCGOZs
51P8yaGKjmfo35fS7P9le136ns/7hWvButB/5Rq/MIZefc9w9HLPZlLOJUxzJsQZ04qnfPC9K3Ny
4rc15tXwYQvlfEDJikbw2pDGjlUFF5XjJSNkpHviMS1eOSlFDwi3ZdKIuDSljbYLJCNuIdkL284q
ynV0ypwcoY1iFdAMBqdg58SUggfbUsfhSLop/jXnQoA4PUiP9Mnaum7gw0L0k0pxLCRJq3XmvLWy
GZUOT0/3za28cxXvyFYfGLm0Gn9+LPg9Y2lqZ+59ARgJ3/drSB42NqmDvSI/6Yryv/jrQNjuE+LE
JJnnPTN4ZH0gfldra7hXb6S1wFMaMVzWvA7rBWaNmmPX+4s73aIZCbnANkS2DedW/UpqBehscTEf
ufzmA3njTIf71khl2DAwDZq9t1jpQVvYo4mcV/jqXi9Uwi0q6qXnvbCEc8IUb45Almgk+1hCodYO
iEWQkUjyPpqG413KJhcdv2EndiSHOTDvsr/l19N4JNp/anF+f5MWmc3HkAqAlTRE09EVwEpz3mBn
4A6AaHBsSpVjOcSQD7wolK7x+BIL/Bmlt+Sglh+uWZq/FoeImq21rhnMWSgUafgpYe1v2Vzb5u/V
x1B3HbrPz3RiMRXaImNVHVkQWfbEzf535mAUw9BVdudf/j4ct2kwJEUAyTuPw/XCeu7wPRTABUlA
OitJZhSq6ufqJyvBTSVjF22b3pKh8qsZYVkDlKL5km3rbhCZP5+zqAAR8e1u1WC0RiW66WqUghgB
O4M4Cqk0ZxYKujl0lCgLYTNIzf5I2TUOVpgsGkAWjpHrlnrd+6OkW1H12ZKx2Ypbn7FSfZFK2cfa
1I7adDueFt0AwuV3qKvInhzEM5VqJNqOncvgWc32OMQE60RF+EZX3RPSbAfZYIIb2cSMERMo1FuA
ymDO2eiafdSG5DgvmsCB6JjwZIkG7tifC0DaCgGf09FtI0Ys0MRHjVpe3GRQAbeHy1A/xrhzmrlu
YDXwsv++vb7VSf/bo0rAOTso46iH+5w7Cgvh2DOFeo2haEVUFwrkozYG+j+2AdUjL1k8JA3uJwYp
TDLXc323YZ8hgtDjaPPQi2l9XZ1lHgghaq6CQJIRrWcAE/9vP+LyBoTHdOgfezrPsyP7CB9bRkzs
z0bIgS9hKecBLswHlG+MlO+FqYSB+wzqQSOP6RLH337NVqHEWk+Xp13XpY8VBU1ft3ZGsS6ez6Tr
+s6KtohPUtQj67iZCQWzTqi7gQz2MmcheEA4v2YzXIriifigNkhSkZDKX56W6aya+fm24N4hV8ER
3K7CpNTfQkdYk8RaFXsya0jJV08WlkxkTMKzExMZ0n9dhIYw1udAcP/n91FmojMBlsA4vWKqLGmI
MlMa/5jn3xPctO4plIR12lKD7yY9JK3Glgub+Hlx08nUwEVlezwfHI4uqE0H0yD9VRcNc+o1rw8Y
1cmFDcNOqk5jyYXAHwMIVXgAhIs2TEU0IlY1lczMeA+zlNhWmtR061qkQEFnHFqWTXCgQysy6ODk
K2RVI9hsE54iMRgJxpF1fs5Trr5MFafFFPRGyK4NSVFzSYdxJj4N+wH6gapFsL5UTDYj3MVN7Mbn
Idc/rGmowd1sPhQ5xi8snuBa0V8wCx2AvqxrfTpE9if3IhDyrM2d8qLnogmdwr40B4Ieucj46pFK
h4iO66BDVJ5ePlCuNVCV+YUxky9aBHUg0EGNfIG64PLi+CV7VYVxEqDJw9ee2nvIBvvzN3sxfH6O
lsMPGTtdfuy/6/L4tSTQF6ZbqZsix53/VoNNxehEzXSQswYOTmL22XDdy9UcbTeYhAHpJiCUTG/E
Ae2IrYGhAKVrMkJL4moGoimwVS7VvnwxbiOfnJXbkD+Rgmr0AoeT0ExxOIiGmbhhSwzm0Cm+OK02
6wO8ARkYPrMI30E8QMGoZ1VBEbPkzW7jHfvOCM8ArYz+v1RAqHs/K/bynVncExQaU0i5rLPkMWTH
ljCIpkHQ2Po0m/jzjvE4eHhaczzk50U7Sdtkg+YZl51kpC5vWXHFYtFJIhx5mQARhL/Rs6Ysc7+N
etwRWyREfIu74+0yEfVSGuYc94xesWtacgfcjCmRuQ0iaxiAkNQsnYwTdBoZew/Rq/sryLt/GHX2
ycm7TVn6OwVb7cO5UvC5F6z9Iigp7G9qi+RMT7VRHy8RlByIZ/ufZ4oDmsEHOtsr4DL4capeZp9g
iPfNXyByUQow/PcjgjTwEKIBuLpDZtsNCQ9eG68pV5ayDc73Da+8xPhYunlkB09xoQrkxOPG0Aoc
oVqoLGVBOP3DFXsIWyBdt6zXsFEGW+AEqIiK2KUYW7VQkJxqTUpWl4SY83vHPuVjD1GjFwCWn5yw
ZSwPwfBMIB/xuRxZn1RLdROPBoLGFQ44xQTtd4gCkqFCzwy2vQnQBwsexqy1cJkI+2Jxx9erT0J7
m6kSWXLzxbEHSlRV49/1c5liurW+KNgKxmcMS4rYroQe/0slqsUlD67Muj4TCdxSB+dHOj6b6QMP
G3gfHTTTXdFzafGer1QQJSjw4bwj8FF/9Z7iuKTa1TiYzkJ3p0BVnwTshic4V3FBq3si+Gv6Jo0m
6IsiN2J99azNifbAIHw0pxCg5rXZz+/tjWxA5vWG1nYEdNm3VFb2GiIfuS6baC+yd5/TsNbm/bgJ
ITE3GS4tEmyQZu3rlOTVwLCxMqPUbl87snXzhRqI1shGPKFgOlwS9OalC8IcEYXDX2hoKFcgeyIx
iEHk7aoR9590NxfoZ6llL0+yXJSfEbaI+0UbO8vYvWywsafDIaphVPtxJ2LPaalHwwLswC8+mKH7
w6ldhYgDtNYZ1vA+6Kz2FJrU0Uxfr4s0c1aVsdKD9hKsJSJvBNqN3msDpN6xPsTT9hBo4Voim/2m
sx2PQ8m2gDpSHTQhOkr3YJrJStvzh0j35OTqUOej9D37FlUSG35/SxyZ2joI+f1+6LnHKWqCLXo7
C40ambuBVmSARUjI6dMk1hV23R6twagghCdrvkVNRNfGbY7jPKo3JEdy/xyg++1Ti8GfDmLViNf2
bWoqamYnc/KH7r7BV5VRAMknumBFW/GhZICI64gKxsAA/HX/l26JeRU1FgmLb47FSNmICVDlLSDw
HeMJzclxuYF8KODgznoxJrk/G7e2hf9e/nARTGiXaPve3/mtol5ykqa0EMwNFZXs2QFn3sAXQ3WC
5C+pqv/k7RuExsaMainoYAVAL1a0YZtkhG7Ob52y7kS94nVOUCULewmQ1n22h/0uDq9vQyawEh0d
cFhGgISCmLYxts1l1cA9ObBR7x0rgjs9j8Cq6vPLQJXxq2AamygLXGoXzFH/kW+n34wIqeTO9Hk5
4efO0W4i2o2kki7XHNWqe0/Te1PG2JTRjTQvU2GQzfkmPEAssHyyi0jjFTJ707qh8aaD3yWWvmUV
5HVkF6uLIJyb5KYncWutiqi/psatSmYsf5iCfGNf6xJiSMCe5pqzMHlJx68GPaF7pWBVcApsAgCR
j3cvv6WoMGRhuuGdiKpmdoxiNGhqefbBUeQ+TsBx2lTNGlB8s3+pD15FO1+Gd1wj0sSNSjOkrZMS
X7o3XEBinyFOYzf5p+0ZiuSKW1yJDOOPkXKXxwxqMCFXQ21i64wvyBa9/vNmGDpXDpzHEgTm8Vlp
02uq6BL/4NqOo9sxwXeKOBjTH5bwV7wDYBmPYQm7KEe+6TkuQoRw5b+KAWIsPwgPq4Rltq92V7wM
fmsRSI0zK8Wj6cCrty4I68c0oIR5pUamSSp8H7ntCclbDT0bH+7eISry4W8q66x5B86N8MR84Sje
pobn5VLIb1DlsPShAVvBILWFh9NdMhFbGxEqv3f0L0rIA3MdT0BQCdpUgN/Zk8mrO/pVjBdbNgCZ
ihg7ufIAcIcKoHSBQ+mc/p8wyrCoNm+7XhJfnc3wIdD/23EF5/KFAYrrBaPgf93VGM8zAUCKIQvk
knNnELlrfMLlWYSpo1pSXgdUfBElRMSgdT+Jl+h49Eok3rrsafUP/gOawY4jzOhgxSxnWHUq5xoZ
nYNshjHuE9xDGzyY+baMbTLPgcnX+9BBxsoPw5WukLYM3Y36AanBGWs4q5Hnjpt8UGxZHZb/9m57
ryJjHsXMso8hPcfjpB6cx4bgCu9NVYexPTiSNhdKyMcWMX0u15gL2MHIn1lHxc6uOOn6cPkYbAyX
9Xx9wRgnB5bDSPFUFtMW5hn0d5rLrMQojrDrV7MRCVXeDGJTbN0PndgPQ8Ig72Vge4BzmxAeWt6S
C1qd0hCTYybXB478bp27KZM3rG35+xwoEbB0lKjOAtt4+dTxpsiILNlmpj7ggb5JynbngsgLv50y
Tp0xHDZJbMH2wmJ/ufJNoV8wKhTbrgzp6mTAV434D5lX/rr5Zobx14uNpgLgD4WULCnKO83GJJ0T
zbWc6EB93LQzCzaElwHr/R2bzAVCAkYIVd+p1IP1MvcsGyXTRJ21W3GurNGn/1ZG4EIH/SxQCgwG
AjcxIzKV4NVkFor3BU/yHWOa3YWmVxk/jqF+OOlFhYUtzR1ccLcW0irx+nd34QgVpgfHW1MXPWs7
Z24VTpQbcNXADp6g8dhJjZ+NCz886X/bFMpuan4zdNt4HnFgSKvtb3G+X0r4xpkeuYQa183CcVEK
5Y+Wv6vbGZNSysJVzUSqsESuIwzmH8SNLgtDASlAfHFxGvmBdb/GHjmK/6yCEbUyOS5dsZxs0QZO
Yy03S1cGOvWhss4F21QaS7MSwInkF8YUSjnn1B71YVchavtZNGcpag9AkCnuQHCQom9DGWietq8y
aCbasah9PfjrKpEDsyhSwj/8uV9ayebBFEgHf9FDHgY4NdCSt5fmobVihs6cUTOg5uORa+PSde1C
F/pSTcN8YdhGvK4ppb5b11/+fHil7bzUUD2W52+17/yqKR6PruQyRZCD0x8IfbBrO9UHOF1I4MLr
Wvn3hXxdSdcm7pyEdxHMCdWjI9w60LcZG6stlNKkRpzlcf0pCUj2E0FDhfyiDhhY4Aqzdz2pCoiI
ZtymiI3QCQM9J8HMgQfYuDm1JRO5YpLf/xDilVca+QUDfifa5guKo7PHzn3oUMHK6NM+kYHWbkt+
+CUgDYGpPm0kacZOG6Jl+vjut8snESW56Uv1/VShwmtAo0g7x4tU3A0ZaL2Vj3c2jgH+V3KAJw1n
XkFquWI/ZMcLzPsmpclVeB+YSjaUcgcgFgJ66gLUrddLVFFoxduTm4jkuedN/x6pPQ9rgxmUlaxP
9rPwTQFHn0S4ldDYVi9rJHpcCHfK3aYMAY3OeLpJdCjlTlH3+cPTiI9kJK7Hrln/rnNOylFoVlsf
O/Z7SkDXWoF5lOFU9ztvFOCJQq3+BTYd2sQB77gjKZb6fqnAkZKJbDwAPsFmNklmk4hDcWMZFpV1
fNOfk3VGIZW8EUPYlIjIzT9E6fGSBgkh9rnrWmqxHA8z6cXNO3hieiGjguy7OdmH4nFOP+UN/CYp
2kluy1sI2iXd4pkSgKDJqfxGgxJjI3Wz6YOVaQwlBQTx/e8+oH3+eK2A8JXmAH7eTlFL9uL4PgJH
FEjtub0eN6Lt+Gk0legEVNVJvFXEdTAOPsg0FqoG32VYl8XZ7017LEhkOywSXyejZSzCuR1yI2fm
aYMlSJv8FMMfJBQDoWQfZTOV6bbgms4c83X9jqutDOJMPWTVvb1JyqohPYNL1xaPEUbLy+086R9O
vQ5H27vPQ4dJZuCIu7SJtL4+yLD5nSu9A6mjV+WB+Z87QN3Cw6TIDjGzufM0b2SWOHc8wMwjDCu3
2hTS14T+y+zPRpIx1jrR5Uw25Tj95q2MtqMKJWvDoYRssmNEFAq5+6fYF41L7YucSMjkVz1/nTCp
zl9t9qgsALMLbdcNL9bCiUTgJI3023plVXxocqzebBmmAPY/OawP24+EPNyGHi4GjXqc0Jf4r/Tb
Yj//NGJutnfrE0BFDUYdoNS19N0xs2i9UTKkBXnsAP9DVFPiinpXYV4mdEYorvXw+BIDefV8iPFj
gOCdkCrhI/Vmh0nAfWY8jnhFh1NoZQSomiAZALvmEWYlGFm7keeGBHkHsQoYaI7CaoTpB+Zuv2Bp
ExJa0d98U2a7AlF4xwHSKfjS8+kdf3AR/RPGv4VNc+PysINGgYYB4U07wk7bPUCV8hEdvd7z52gl
dNDDxG4gxGxZJ4LQzFCKJoXv4KWV9vw62WCs9jm7Mtxz/YjMZ2CGLHvN+x6AO7laZgkhvzGN1ami
W4blM2O9VvmtyGhP6eCy8ANROoHho0mC5SIwPPChNvj2e0+5Z4NcvKbNX0P8pBtVus3YztnX3AY0
7XTLyrM6p//uv/pg2VdiHRcnw8giUiQFuor7LQxFqWX5ykd0pUx+MZEn7dhEH0d/jtps257Ep4TF
59iIFJ/DvH2S6QxOrrsn6RXvLjVebj6VoE9dD4NJCouV0XJMfwCIgiM5UuKNAwNs5Qkq/Ih7xYJo
Le34Mvr5yiPF154ulLCOiNB78cxqhZGkAk6Kk0+Umx7ElmcfwNxg0Fd6NBaffHA6V5lC/DXjzEO6
RJwQuELNwVgOoWjV2/+xOEtAlYVEEftkxXHoJIuMS9KlpJljLL2F8CCIMAtyANWDq+FYZYPgj3ie
d1HDHoYnADmu0V00zDShzf5UwaCmxyScCFkkOVneS69RNsgE6P0w+ZnVA6RinVlzMNP8vrIQZ7Wf
JfDoL+6tuq9ryKqfHFcTg9MfBxuuF/kYdgvL9K0drWTdBEauh5oIXJvjDGW8CCyA49++xfIX6wwt
doDTVb0ew6D07GsSNMiCGvqzuFV35UbJfU91Ayvnm7zs5NO6KleoMlh4cHvaR1MYWFBZvurnbdWh
mYdqP/DUQ99gaDTnwfiYQfdLHk5VugMx0lPB5kTHwvFSlTJMVCjjA7b7sc8s/Dc4kN0HA0VE937d
/4AatvQ9bzE82ZhFi9dYJBkboEST7vpdKzA/vSFOGDcSNdtLnU2PF5k/Vg3QBEMzFFy97o+0CzNV
NIJA5VY3sy27hWU3R21osqAMbBeq2Af91v+/IFNEQcdT8r2NCk4W0bzdC/EBRpBriXD3DmJEZaJD
PNa9zB158YVEOb+M2ErfxbKDutujfC3UdMSy9pjofWKwKveO3aRvnfT6NmqZSMQLnC9DnGZ8Xn+M
doaJP16hhPrq9K9PDvFVvdr8j5FZhelQMSqHOk6mfrHEYaYHDV2NrUAUA1tZy8aPPRD54f696TZr
abin0v66Nq7hhUFGBkv5FkRhypESNnWD5EZDPtOjxQeIyJ4CqHh+5v0KdPEDtLHxw/Rt9SVBPCcB
xulPkS6Ov4j8e8/H1N78wKClLu2/0jfH01BBDaT57QHWEyAGGAdMJvg8f8AfLqQ76kLKOcowjFYC
LZXVzPhyY4Cuv1NWJCQ3ulVzIFc1+8Yw9ax4hNNfAyS8VVwaYc0MLZA37szQVSXDW03yND9cWrNm
Jfk3y7K+w2pv+jjZDPAYOy7EgLptNAbN87xxbXS/SkNZdujwxWnvOScRXA47MekZrczAYy5T1Yu1
meEsJyPVvjh7ELrWHCkirqD1VeU8prQ57qjLDbiMScuf6iY5+2bRYK/dsVMr6v59rGjboddElMWI
Kd9ep3iKaWUAiQpDLHPC7wTTpdAEuBnw5HGQFJLXSelMml2sShVTH9Dg2EjwOVj0X0VsTB9DhYIy
qlXEwIeeGuATDxgGBN+acCjzpyF/cHyqxlOplAa7Br12zsqE0UjWXOczh/geceeF1Vy4aKjVNF1l
cKSUQGWXJ/0xhVnhMFX4PQf6EboIU4AXkQYZtFoI3xn1VtmnWxllKRIBNTSNO2q57c00t7WgwcfG
c+Md3ntMQkr7fQn282TZmG9KOBSoTdkld5I8F6t5mwV2uYqVSjQA11zqiq0KiZJbZFWyfXs9qzjF
6XBfKx4PgDXm0/ALjIazsDOoXy1PCTx6VwKNdUEs4LgKq8yqbzE34oTaB8q1kD6VBOgKz3CAkdFC
x1NBT//J1t7YyeMgVvu6dif4MAWZ/7QLBy5WeMM5uU0PbsnLF3h6sGjsIx3npXAtw9OlVcKF6dkP
EC2JcBGB6w750o/Lc3zXZ0+vFMOsIPsKMMNLBCGJWwElnnA4xvufgqoX7Z9uSnS3damZPuG3ZHUQ
Adbl5KiY5GKbq7DfFe/UDjkmba9yssZ9Q3AqLIczOLlHrqy7KhQ+EnKMWz4gIHDyP60aYRR/5ya3
XY1JGDYP6I2S1FqEVRuidDoyIQbqEyVXNxJe/LM5OHwIRbGdTeV0m3jTfkP5o7OUyJhNgIhKB3gT
t72ux3sapBTpPkopkfWE1RIGyd6DzuuBnw+E7EWhTAmNpM0c2dwsJ8CoJcrO89IDJJbOh8YzhL0C
d86L8F6661WN85L+lncVwtujelvMSeKlUZF6QxFMdwKhZrTJW9nuPe8bvaUZ/V+3D8N4bdznsfrU
9pSLRaLUD0lNOtapTNqUb5WfY1xqXSZa+lxwkDkptaMCQBnKC4nLHOqKqhc1rphA1wpHhDxlQ1pb
b4ZaF5j15M7wsnrZNERbVGqNvVM7Pk7FHrTMbD5OY3HwkShWDZDxVpxemi6Fec5dElbmlA2F0Vc3
PI3tZiTdiE5BLCOSLxCirWlF8o30bAI11ODhwEsnAfAJNVElRb8hTo1YQ1OswmGlTuLE4gZb16Jn
DSPTIqAoFfVcMGPfh29WzxSn08L3TF/dHU3eCplxFNU99qB/wZQgzNuDW76Lpb2b2wuGa6aIAsJT
4AIH+7opb6bfHuUi5U1N+dJJFY1Os1ouaiSjcaNrEiSD3IEr4nA98QogZdb9igkltjeTnOwR0Wnu
Gcdwr2jQOx7EzlexQgpTuobY8eK0/kajits0an0mp1YxX9BqENx1WozFcXJNCVh90z7XXXXyyNE5
JwQcEvSlRg9lTM2IF2Xw9rvKYM5Z4JWDjWe9R6kuH/fpEngXdPitM+t5Kqm+accVaEu2Cdzy1f9t
FAbCUCcLfTP73hBYedQG5S2Vdewk6sr0EHyzDyBCb3naMc+n7SZLfvF1leJgllwcgSA4JkEPGtuR
mzidnkgH7wWYm09A9v1Ia1tM+yRDK+Gl940g//di0WLA9ySxA/STf2J6/R5Mx07g+2wA/uxbxYpN
Jt0KtHjwQT/q7UDGkSUJ2rBLqsiAiL/rmNGCjF/lhM8Ryo7jFr7WJrqvM30gq18C8PM0d3loWJ+E
mO2uZeO5n8v9RH51IYi1g/WAq5PGTZuHEvhWcQwYFGCTijcyENdJsRAos0R6udtcUng4iS9wTFxv
1OSBq+r5ROMbOn4F6bbKsJMyKhXe9yYqCW2sGFYgxz7jadLS/5Zrk1MxsiyjLtAwWt/7kv5kGO8h
t0iuCrED4gxOl75/mkYbJiUQH7T6v8r79kCuTQXsPrPg4m34OO5Z5yvZf1WdwJJrjfOht3kDeuoV
QQ8uZbKLDdwje98yQuAkgQuoiu8YhvtP3TH4fvBu1cCEtJfdmvTh0XEI3ACw/bCxs/bxgOgZIj57
URYzg9EdlrghMEqttWi5gE/sOz6z6fETGdV7AGlkcB06i4TjG5nxHuShBiF8nCZHHjNtruPWFsO7
GCubZPRT0LM36JlhoKo6eJVkEnP+uOyJc//slaZG7ESiWXl6VYHf8y0iDZLkF6oqyxMvoQUsMttd
TFqEzjT212s3KG2Pcrd1h2B5GsDPrLSJPJz8KozMwwCT32c9DwQq9xsEhGQx06d6zFLITMbEbTVN
7F9NeSRN7zAPmAi2gib/NXq7RhtyUiypEzbm1BcxKrpGRSUiD8SxNjNITwfQcFfNlzXmlr60Te94
SzZzZokc910bQ4q1KNDPgxUCrHnaZiVM85PdU3s7blbhBSoVyuNCI3b0yAfQ68RJdl3TM5oMJsci
YzFHR7QuV37Ynf3hOGi0RBvXYMBxsmGNHrjjGAw+n1GeMUjNB44xcljnQH7E8n/09sM+dhlsE0ph
5RJbjYPlPgRCPEUPTobHGBUJa3b6jiCbScKap4b6yKqZPqYvy73BBCGKMsjnwEO1qGbAXoR6bZH4
TVQ7cvlC9tTH3j80MFSEr3765aCTi4CU1LPLL4uDuvPmLASr/ipiqfU7i6VV1kgRvvbFCrf6u5UH
pzh26O1OsJ8vjszRBa8fAGJ9U8jdvDpQsPI+achHf27E+QldufIbi6G7ZMD3x/9ZrDsER0MEqQol
YeHWziuI4Fl/2DwkBAIsW/ohGcpgPcjBbwedk0sOkRrXWID/dnqTtrquW2DrRM13Agoy+Dgima/j
+IZFBRkHuIoQqvEurrTWEWBU1MaSeQ0bBDB7AGkOp+C39vvcDp5bTvNyooMf2sCAciVMKelexVzu
eWDNvatclXV9nGxYSn3R3A67V7UXCH5RguXDUq3SMlmCx4ENVzAMSWA9Jp3kAc+NfGA5M2YMvo7Y
8Y1suSoI+d4mPAyd6qcoZgRVTU6ckDknmCOkVJXf9sfXhQ+Iwz8Eku3rBoLHVNIh8EGFKKcOPv3O
eMiFXbGaz2lOnV5CAJtElnOxqTKD8pWWcNy8bzMemcuYCvjeRIRobn2MuWpZMcrFkaJz4A4EJmkG
SHn+A5NwCGttTmbv3vinptJpfOD2gvb2LXrc4YHFXk642FTVbvBy/OacNfoddHOY9tRyH8O66KUD
hAuFHKIa4cWi8Naa9H6qHDvlEW6B6T+TFgSj2fDrVmEC9bzepedw86DAjlQ5tWIasfsAXf90BHvB
RqrO0ttVplD4FtqNqKDB3MpiH/lXeOdDfwa1gUDJ7l/nU8XxlJwfiVlroxrjXkwsk7fzyZ2zj6we
Iu2x4WUIElc8l6iXzuFNyZ3tAHsXVib5VRkOFqz3/MMWInAizVoTPeO63Le858ZomwZQwRCUo/nJ
K5k3RnSgrv8h5ev+aOehzlgZI9fgQvtfQG94xEd8yMEU//cFT9AjbS0mSGKcC3RQieMTLJ6TvEn3
sRfKkcFTUEI65a8U8wIIO81ilTPUtrFpkXlFe0Lqz/097gpH11VN3+ajZGb8wzL4GOQQdAKft3/Y
JqoGV8LcZXEb+tAYR3+mxMQjtSh/Sb9D3g6ifUaVnzfCHbnneLcKvPydR/kaTiPWDXQsVehC/yoi
rA6eBWGQuKerv06iv5+v1gI1OlKXertB1vo+ubkQI4orhdXi+ZALl+hpHqDz1zh6HfZr4JHhRX/H
fsVbpYnuL8EpU0i8auvfL9MWa7+b62ihcfUZU08W9jD7Elf2VS45nBp54igj9zl2IziZRfSSBGxK
a6uOurkktwFStO8KDoVnY/+Q0cHymauEckgjU33iPnyd1lou/T6DvQgavAsRfXM3Luv8WSBypKfo
XD+8jKXYpIxf5mckR1ce7H3CKYH47smIMbHOq3bRLGXslLcDx8dkeg0U0JI5uOy47lVNSr1syWL6
T3l/FhmG35HfIcT4g+Dr+ACGfl3kFC0s5lPlxEgdBQEs7EdBsfTZRgt77VzEnYPrMulPizYqkrFn
2FJrIQVVf8zumDapoAMmcsIgLgz5oz6Yawt6Y9A6gV6fQWlzopV4J4LIC7NJP8DI3P2Y7qxn8NPN
VpP4EzMfkRlbe+VZqO/6KzD057nYPsN3H76s9eEOJMbm7XqOj3hQmdQ6gur9SKFYu4MNkBJ0yz9C
rt81HDHqtrkBUXwM2t8CyPec+NOyZf4K4KDTjk0sLTxQCPfHsEvhZOYT4xNDSkDL7ul4KnuECHw7
WOgf0R338TdFnNpzKejzeIzUW9/zDz0uSGhtos0eqRqBpp5h/9RX0aFXdIZ8JdDn1MLppICsLum9
KDwOAirynTFpn+LoHjYhKB9n59gzhVX5eQ05DpT7i4w+6Hu+lTh7BywZFNuVg/0TQo9FMT1yptun
4yrzdxpZSKXYs94djyVv3Mb/3C5ebynXeJqDYR/5NLyJJqPWZR1XeMR6tClqoeqFnlZPgnuxslUO
sjhDFbpq9+6qRGvJLzxPW8ePYfjMEMeoFlDm6rh01dQcccjUDdEpgLMrlObZioCVy9JyQ+Pfdo+C
n8VXTuRsRLUL6vvL4bd+/A5NHdx5V/89KWiGq+fKNGyN48d4yVda7NyCHAyDh5fcSrE8rSSy9tmH
ejNnXn/EXiMJvSKVldAQgui07IgqQrcgNHup317XS0PuZfpBoay1ryPppwq+j10nmvZclfrEQI3+
cqWQj+25EWjgxWGCY1x1xG5chVwkIyDneQx4HwcVfZ298S/sHQHpnLuF16vYVMcNtV6Hd5SZJ34h
QZnFVpQdLi8I08rl68o64MRNPODAHek1L9r5Ga4uv4xDn03EaLIpnPznLSF23IibCq85tqULV5ZW
ZWLVAMhpT6Mr8CjKGEEngEIds8XqQfK4hjD+RkknbbzBKf1okBvcZLOXsA6grQLIPeKSw32Cr+jy
7vTi6Jr2vWHc55wF1RXWxN5H5nyGi8VRvnVmd5jCPKaQCBr9HVPmzAv3igK0wECVWKPUv83NlYFo
WQg3+H5MXgWihoJBpplZoEEu0xzyaGGXUyV0reTCk42Cothv2XCcdOdjQAZGbzzfMpnZIhNMTVjE
p2VTUT5mNj17DGVRw+EORiq512C5KhGDlf6SC3ndH4Q3BHeMJ9xeyOTBuMsmxO1WJ6VqYIpT5GNq
+yFPSvYv67XBR1Ljs5dgih3z/rBTVfV9KFywLy0hdEyGjJNtpbjajqccoiScfoFGKD9eiPbSSvfL
iMg2GzNkblTqrD5okCyISuHEMMAzpibQUn1MZYoC2jibWIbSowI7E7Ik1St0wEEq3WkCpc6norOy
eZXo/+zY2hYp6O5vGr7xVq6We1528IwP2inp3cfzTfINaWQFWUbM6iAt4UEhpW+tPMbTR6r6aDMy
W2Cwj9KIM8PLCfjb2cxS3Xt5woK/Xy0wbgKo2KJN1Cxnkq0XwvEpBSN9lUUJGSnQ7Zme6ixYpc8q
ajthSBFvXDnxvMfVoT1AX8CDqpWJayPu1xZbKErJK4+mTVW8WhHJ2csKs0pxvbYgC8za2EsVmM3M
8/pumY7Kv6QAVG09Rwd8vgvq3HCGAs/UTpX0gjUDnZHwRr4J0TjEcdui9OAu4vUl6SZHfqVyYhTV
iyLzMP3V11nNp9qOhCPjrcCqOBNoUl9CaF3HtOONM/4GJycmA/+lp298Bz83b2p0GeBtj+N6kUis
VKb3h3el+jwhqHMnhVLhS9lsv2QtdsTzFVf22Bx3UENFtTnOkOE6IbVdV//3NCyGdHCIzRy5oHPD
52z/FPh87lkT389fzpKTQvdxCylwzBe9vDFl/NgFSejMOmYnOJuqKEEGxCMp8DfnyI29ivQNyFT5
o9t09lL5zBekt/dXI5KHRBuG19zAc6wpXY4Qab9Z3pjA78YF/z9FlJnqdP1A9E5+tvrCyPu5bDK6
U7CcTsXDiT6OG6JbH6pJXYtT8oR6YXjSDdst7pUdKTVmAfSSBr3AQdmOXhmjYnz0APj4+pITkikC
tLGXidVIppykm7nEwpHzgOUaHAGwqBEk+KruNwGAYYKJ2VFEIAO8sEgmX/9nghrYJa7gzdkHo25/
ilO7rCNUmZeyTUUkDRpS2uc+USRjVhmwFzIOFVGusGhqYH/pprXD+sr8WZtd2sQ8eHf/sZubz3Zu
hCysGdwXUhlNQpZyQcS4DMi78vcmtufC9sVOd97xJNqZICHYJttEM3zPOGDdazwuHPJYLMQosnYZ
MVzmjxeKNUVO++2tgSjWVdsJ5K1clAASPkQVg7/Mq6wjjfksa8zFZoqik8eLVFZig/kkzEpQb1UT
DCDTHGKl+CWVpQCL+yWXhp9eOctL8tWdoG3rnlbbo0UxcnIr0LOGNXmyrksGtVbnHmsh5wEuSomR
8IjooBQcOzVMlMHx1oJrLf6oZXQygjXUFTvwp583rBpXzoGrFZqxUzK5UeX9+R2L0aZtQMqmqsdh
2QBO3QkYGEd5KlHMXh5s1gAhrCaG3mmjzWLmFhFih6BCLAQN5A0H2GaEq9HX1hWn5MS5VTlR+PuR
r2f337guqDF2QemwfESVN8EIfhA3TaToXgk4HqifXAXBdbIbXGVVSkwAQHMzMKayzQ33wp7i5O8s
oB+X4uq3pzUVno1zNhC2JPTkDR2HL5tLW0/q24+HY//Ux57M2vPsgY5zWgINWuldnkOHj9gYbxIF
pzSr6Y3G6N9vgKAheVJbvCzfJgNmLIFfmqd4hy5rzO4T4BG2rxytZZ2SIVro1vwLjQr7gxyBkA8a
oB7+I6OJsFP8ta2q7B9tgspYqYBTkuhd+be3V47iImIoatB/+JDmP+jdKZeb72cjEBo8OCPTcefH
J+P1Un1GfH1WjYMhg3IjN3wWkOy4go0nl5y+lq5I+fv+ql6JvDfcVjC/HZ2T7nPh2uZTQDnUnQbW
i0Uj/6dbtYQbp7f+mp7v9ybDtH2IASiuPM2Wlmf4NdINJ87bxfnv3usoRiohjTfXYZ/8IoRr3Jer
2Gzj6smfGofAjsKxJTEACR3Cj5bnk7VnUREKoTYOf6aANvjvKO2df25nERBnpQ0eHACuG7yxa2fs
kdg71SH0GD62hvs3SjqnxosAhbIrkcde3P52KOyaTaAYD4uqS6nHuFAJbZFKXGTIEWwscYFdqaGt
SZaZE6nwEqt9AhTybSMk1RosAeYM0ZLSdmrVEROoTcNEl3a3GB4xWa/u9rfB9mUMbR9LrllFdVGD
nMH3n/FVXq0nPprKoilG9KryIXNk61eswQSg5eKr1E+1BifUHNd7SIaZSHj9xzuU193QR4l343GG
Ny1rykF4PeE2drHBTDLM/w4RqzIc2jyou1Usl8XKBxkZHTX7exb27kDM8fLqCVAQVLVealF7j0HG
c/S8ZyOJ7P5vB0x767AMy5voc3mHUTQT1PtLtqFShVAi3Jg0Hc1mqAUojm3AbI/Zh0P7sBIe5B6P
8rF2fCiW35DvUft8G7Cz4GJ5npW4L2sjs1QbXxF0wfbZ2SjniTlGVnuJOFwYJuYu49LDM6OwiJ9x
C0RnxrG9MtIp+LgmuJpBrk5xHAw7Yv5GSj9K30DPzvmAMeg7Ji+PeeUDEhcH2hh9G3pLaaOqI3O/
JVF7XfelBhEqouo2MEuQNB93kdgV0WKRPUXeYY/jozURgGvXZWS13YmQ6rNNTua7Z6l/H4cYjfne
bFq/nQpLHeLrMtsGWquczxNEnqOmiHsg8MYDiwu+PpTB3ZA8+KqANm5dcQR0//YQqbjP2Z9U0vax
ZHOg/KVwkP71B8pHdj1KJafuS+d6sYgFjN5nNYCUuhaawQJx3fCcSZxGakOEDsSDfa8IPZxsZrI7
fZBKY9Bnt+rcXgNUelhYWdyNoVJ3uTa/HvHP5kE5+MVMSk9H/YZuQOVNbfQ+hoAav9Cdoxeg0yCJ
g/xFykdjNcYSzsKljPQeqbXizPwmR4PGf3ksApcIqX2UinYSe8Wj3H8o+ZHHrR3f1T7fuJe3/u01
s590kCc5X3HTJIlif03L/VA0iDnCHVDpsDFb03iUVHeCInT4gWPmLdWry+QcYcny+AiiH6Z/R6Jj
WrmBEyFW4AyIy7jKUa/arn/pFOWgO7eFAlW92XRTJKf99JtHBM2O81l+uv7uIsKcR+PxeMuePxh2
m346kkC5g2ecOivb8zp59hsY7sM2BB4OTOQVw06X0e1yrk0qArCeuaCGL0nFu+9cDFKcJAuwMeHJ
GHlpwkXYiduYd/qgnD6f9/bWHNQg5lSchujtwrkflzu8KkXwvY8ba/ECIb3SQiyMuqhJIXUgPWgO
d3wTtTSjeMt3pSHjjK5kB8iUkE9XKTSuFvsr4RjeNlRLFt/th+phyvvXsui4qN53K02g0mYSV7X6
GQ0GTwuJ+m5Mc9WfuhJANodAP+QdO8c3NqR7UbQ/kgDBTINuhcScrfih6c/ddHvfjfjJUspvhJ0w
l+H/AP9OMsWBpUQABrJz8Z4l443+Q7DCSzpukAW/nn6oDS/7L7RxTTSSpUH0VZ83/BWTR3McmGiY
Is12N1+9MNeukYH9czjzy1fHeGGEG7aBIyQxqfPX+tQEGQCec4Ww333OURLYusbU8IRtc/OWO1u0
TAktLm/4Azqo5xBfetD1/f4dZHza2td0DEsa4R2TcThTbcmwd+WdkRWkz0h0JMs8u8p8Vdn09Uq7
rnl4ku4x26+tw87OjbEk9rXo9lmA4x97b4xIFhH1QtTZeIdXYq57Uq9rlaaOOpfsxGuKVih0ybRN
hB3m6y67xe3pYeSzstPXg3qM+oEhRVDCsMKOoRSkiE2HLCVM0DTVHWFKhohGSyNnRpQdffL+/Rfx
ug0IROzoZYj5HM9DhQcLHP4dtz+T6fdZbmb/L47/xaHarVvnyG0eRUPacqav8J8WFP6ttwnTVT/A
hCYlgpsKsGONTd56GvYEXVRak9xCTzRYxr8MluT1yvzea0Ai+XuHAmXGTCyzpAYzAR7pRh+4XgrZ
GmFJ8mHYItLuAY7Qke4VINJ72kwSNWZdceyclaQOHTKrYvyr+lVXel1R0epvn43smsWY6+TMfpj7
b/eA85NLQ2i3mwq2N8TpifdN3aa5Qhvr8El69Q+MO23a1sEaVwgcRS5wEv+xpjDO2ljoS45ydqgB
oaN2cg5rQQcoHna/OtxucJHEvI64ydXTHJ8l462rnrjuSGhQqwbrrGx61SDDjGpmzJ2d+uDg7MfX
HXmq09a3po4obA65IQ3vzHDRsjpNOxqTVmSehf+ij9ZVYmjshwVcvhaFaNTOZxCLRmoDsgZUuF+j
vNqyJNaL3T/tk0P0gkkSSfsRaiUD+YrrraQ9qExtoUoKNGhwOToXCkGbrWtqjtTFhLkzX0ZXTyI+
KdymbhILR9SojhERKxEDuMzVyxP+Xn1hT/kzUg6frTwQcpfFzzky0GypXAWPTn+VABVwUH/ggabM
UHTEAkmPSHh87sbcQMiczZI883k+L67vp+s3P6JHKVpAuJyg5uP9uZhXcGzvPnrEf7Eox0QQtp8N
rQDU7B0HovJq/Cliun2QRFMJ9IbB9Xoi51pNFKiti4saBNjzytmDN+M7EioZZYVqmI5EOoMEk9kj
nzPmNQC1rpluOGWdjsksEr7nl3OXND2Ft+hu6vtvVLJCpflonDyn88xEfZF/r1IyxOeU4vD6yS18
aW0aEcZBhSk5/jFteIF5cBIHuD/0wdXE4Q+fEWdFcPMlQmmGINZuXU4zvr3pc7vugh3/plmZGCw2
hPlBOvdIcAClyks3ou70NYxLU4Oy9OM4EFtVmUCUi6WnSS4xbO3X81CNk3CcwNb70/Y5c4eSHI7o
hLVqE/CIsw8iZKO9n0GWwNWgZ6mgheEltCv9IBaMEmEjwFtIqkG4XzBIWEy9G+peYDG/h+Ww0MBZ
tSCWIbAgq7c9y+q71EhT0jVnztgX/zV3CvlJrB9MdMDScxFyTDneYxDkZb/BDgNFlZbBnNUzCXoU
By9Lmo9CJncDr0rzrAeOxDU7fkur0+UF4TVk/+xHCZPo7O0uIFv6tRtaDFGbKFK483iUaqeN6d0i
i7cBdVMBXNCzDzDhcPUFDvxxYy0Oxt4fRfd2ZQPX61dI0Di/Ct57YVJYvEiFuZKAtbzz5rZrTIeR
TS5AvMqTdDbbaa4O+ls3lMOT+uu2KCoq1bDVCTNj4n1UshW0w+9rE4SDOxD77hmi6DN9NuWYJ2fF
qupQQgyd7dUZdAheLxTy/U66NDwk1AEXMpiE/ormGcfbm2OaqaEUo2matpU1lpxsqj8QP6I3trZH
NJUi5h8sR8SNLMAH4XTD7W/52Wvmno/EcbGepn5w3STGfbubtqZWssC1rOdtaeYWbkFo1KY67t7o
OuxYPdB05WnveTXktaLnsgbbtk7Xijfg2QWDHc2/M+c8/0R8MxP6ACNQlgxb2PNvAl9Rx28s4Vog
d2lZyPVDAOSiTNx87g/UFF8ossZePLFWk2wOX8djEC+mkTv3xkYIdLmik//D2a/v8GZKOqbpWq7M
+/5aNFW5JJU+vUQycCf4hvQQg54vnSVH9J2RXyNCHL/SeHlZ3GrsRag86nH+exKVao15X4JL42Ck
mom1PTTd7IOHcm2kzjjbjK9JNrmDDipxA6SWTgz7xx6Y+FTcGRf/8Ekrwlt+BDSkBkwOVOtmfYdO
pjXuNTpVvBPPaRcCShLqhlgnphtfnVYqNJP8LdpK8zVOOfAXCVKISCZXWeFvUZLWk2ZQAB+56DO6
ICikgpaslBaLyTscDWg3cseRhqMTI+ZAjLuSG18eSRRddlHhH7bhbd+/Vq5HCyZdJvooQJzIcNSI
pRgfV1IAhRvgGMQFKcG3t98NIHY+wyzGMd9IL17SSwTw5DgyCCG0w3pZBDctRwDw7SIRT4p7wfB+
VPCcgaigmqvij6FEqqxneLELCPK5ZGIIIjktEWAyQWIaxqqqk1QpyLWC7ubOq9RY1XVLD/RGSEEA
n1VeF89msMjTU3cRGcL0QjQt8di5/1SUyX83PKEuK/LMqHHO4yKaas5u6XSiBnA3R9tnJWALytPG
SscUYAxkf4lKvlNh8ahGcfJUe2TLujMThKNy4M4sYO4zyM3a4eAzNXb3WeQ5+PfyNhQCOk9yv4yh
ywGAV/TSXvAo/Mf+x43wt+99pGFGIylHbcAQUqKMv81z4rfVojb1IN4+3BBIrb2WP+4koq801tY3
WAaeBTMEtA1MQm+42Eo3dN58fq7dS32YscnFLlLkEpvMICmmx+NrJpQdDsmfz4oUNVVn5yImUQHi
WZqUQsRy/8Dnah2VggY/cfuMIQmek0X4HcC8TYppQJljzU/Yy0LqNa0j/WCj/kqobmx/XeX+eYMw
GQGZbNZWX1ca+Vv6U5km184ar0mUCQyHlq1TOp5pvLyqvV38ryIpxWi2bhp5soZDINDVd5LpurF2
qh3o8G4pTOMBp5x8TJeRTswwss6uu6AgU68xBq9/BOWjeQq5cmkxDyT8aWrFvl5uj2eDNv3K4DIJ
iylJ9V28psHeC66oQSBRhpBcIfFv0tMaq/VJZWSPayfiTjAOClVy/ef07n6AF5agQaWeMS4jbI8q
r6+B2AGbGrniiCvTedWf1lUFui1sNJ3MVAMhrE1m3Otaykq7zsbii9pee2FDDHeH3EQhbPqVQaVI
MRty/fZV+7TM0bHyWAcsMhYNcPvm5WtCjyXI4EYXPAtYFPyLzx5kNnuJ3f/8Qttx9fGs5/TSzWc3
meP4J6xSu9MmKZxXHNDag6zHiG6FDDm4pNI0MGgrCLw/1FZZqENRAAQPMMc8EvzJnqED7l+a0ETS
4Ov3dEZabAHZi+v5oIeiv9hyoa90EbFnmE3L7M1Xy/QtF2h1aSTCtyV+q+rkvB/x+6asB8uKfL4b
Qs1W8YJo7MVyNc1fEer+rMIuhJVjdL5jOvbkNaZxjwM9CeEtPJb3Dj4+LvdsVy4rgsOpgxJq7YJ/
236579N4RO2+xJsFGrziUjOD9UaGughz34E4S61G13w71S4Dot8Z+FVKCwCgcvek/RVRJk8NF581
/8RAjudNUWQjSY/cNmUmUuKlmuku2SDz8D6CHDMg5JMXFda5keexvqhztbnUZYMKfas5xe4LC9zi
EPVRLl+B7Wse8waTJJNxnNxk77PvbjIlbgSgUaawTeepKsPoZKCQmZrPBcKl2ToqPAX5b91rE9KY
YZi+eIU7mmEQ1PXJcvqsg9FsYlN3Xwz2nKJ3O28Th0pri1uE2hyuBmnhuPioZY1Z4eMNvhd+s/PH
uYkLdgsY+YUdCTjQGtymO0UYWXjRA14MpstdyEHNDn2xUzSW3Tb3sG3ZHbhZ8SzPqgWBaHCdgTXB
T6iOM2FZduGtadr0QRRxF5ktQE0AfaRd99nS6orZj8B0VnL+eZ1qL4JWKxyc7qfmwwWu+nW7ahhB
M6G4JrZJMzSxzu1l62NJ7RFqsaS3HUWEt2MB/jzShhV5/JQ+7Vkm5g21Eaq+3W766kfBo8AAWRA2
ELSvMCqrUBPCIEmRtHfuhMJaE6owRyFuyyk1t2hfj3RV+OS/Kjk7AAY2TNIPmgmkPqGGLO2seh9C
152v8T+RXmUT1FvxZ+/qqyE2F9H9vBctWCs/nYuNXPbm1G+xVHiX/F7Vg91vNX+gnufoWwhkMWcg
J8U8XTeDO3czQC975hU5kQccBho82eryTSk28RFdgVYQb38rjI+ELmeNhW/FWorJKbg56EKEuonG
sNTUPqGpviIQXAIUc87ff37RFn9lMvNJUYmaUHxyhCXcZxJ6yhslbolLTSTeoPBe8lBPcOmoO+tc
5XUFqGsyfGP07lFwEtvVeOsFOqYC+bYFhKb6rdf6KApP4TRbs0amqhfGvpywVCmgOo0LP5n1t9ow
cOckJxl3gPfVFWHOv0zoF2WXGEq3CAskBYh5d+xVevfINhFXwolJsB4nETCiAgasSIrsba0mg3LR
6pOUDZiH1HG/HGJCtLGLMVCFhDUuKL9otUhb8RTzza41UmkNXSA7mVP0nqiJ2PE4vsbbCHKiBPgP
8S4wHrF+WbhBJTkoqxjdgdpFmwqNdKDAkxj7I2Gh/eH2CexN6E2yYPCY7pRXOOZ2DZcatno6r/8G
sglFeV9e2ZtniAaDmVww3NloC8O3mTi2rYBwLt5If+BxmS7O1eDriiz9CphyjRiaXY7mIa7BRrxO
MOUJ3VH4XPcRoFTTFRiZ5/2MKgUGYtjSa6FoVITCpI0s4m31s8vXhyv8T3Uq7Q83BH37FT6mbOX+
pQgyTVmbwmHVO0I4EzPXboSMWyjgSy7I1T8anxfceIHeNsM2RKDsKfGVd01G68uiwZapCZStPOQs
1LQGddTbYwns9z9JedDi3GKWokk+5zMcTE8H8ahQ4UeIVzBK+p/gLD1F+vM7GTkfbekYNEXWHE3K
x9e5j58mXpPIw1sJWlaP5KRaWh0fApn5OdA2y8coZMonfjmgkBUEg0/sM1+ya80tGzGMccpc6NNe
yIX4X/gY1TQYe56i189i4cnG/HX92epBiqDJsDta2Xc9IwoQMySunyg6KoNMqC61f81q0nTdum4F
BqsNTNdEMPe/DnpTpCckzMOdteUmrS4mRrJh/WQxOAK1V4ZPMmcSsA3vhmpYAToZ8XNV0PCxGzPN
BivBZ7FfqYDFamU7hnCLFurJSMCZKwlhyKFnMhNeJsFNhm1bTswr0VJ1bTVY1VpcZVLoHju1OsIf
LCNg+6ljbMgczECZo9AVNv/OFK1Jlhysb5OL+zVtA/EEEeTShKHjNqqEHqnDEFpeRDMdDjcPhclG
5NZUZOu7IXgG2NHEswr6Lz3QFwabGGrZjGZiRHHic2rfRjE2S1G+BDSmxbY6smlUT5p+fzhhmJyz
OhhRqGclqwOo1H6fUpIfusaO7i32N4+X3rXOBqvwtD6nfZY930RCf5PZapMGXMj9foL73t+qHBBM
Sdv2YO7pT6R2Yd558BnGcr29E0ARefsd/vJcfWswGJhHidR4rwMtoElA3RAGUYL4IICMWI+IF80s
mp4aNJABw5Ipg0CWtQkUIMQ6PmwP1MeG6YBZS93msv/2PYf0gh2PvYHzjXl7OEmiLPV90fhmRSg4
DzwHpox+HlAqwm/r7HpR6iXVebs9Ac5+mkiEMNesuLwFOCMs2HrHaEC8VehVQAaAIJj/3R6SwIFm
5CLf9JuPcSzz7uLab2GELSl66+kk6GhOeyHb8yzqNRpvQ9PaVT0wXzZl/UmysaHj1wUQEKEkmb5U
8e/hiM7Hn/2dzdw9PMbLfoOGflkH86t7CVhf0hRTArO6YP2QoGZgemEvaM+PDnxzX+MsZBOJ5tNX
02ePLDJZiBygiJkAUnEbEzwsexAL6Nq8l8aVmVbxZ7oCvNvu5N+n4nNiMo118kLr3z0Tha49c/Ty
IM5x7fMuGjz9tlfxbkjD7v8l5TQifi2twPmbDdfIIiY5C4mlwRfQR4O+PWR2edknYN3HoNCdt237
Msssof5Haeo+Rn5nDcb369wSdVdj8xAdg3AT8LTvY2llVk4hHGohFzyPT6lXuHL46d9C8/UwzOkB
4c1hnq1uHj3t9lfJ77c5O4j6pCb386Bo7ijzyCNu+bOi3ys4wiSokc+z6HobD4ForX0dx3Lpt5XQ
M4+3Pt7otdyiKP+MMDLZCoiTbGkwKrJz+bCSdt3xCmxDKSt4MYJ+CVEoSaYBMmhthodKKOUbQOoF
tVDl2UrEbt1+kDf5ijF9Tm4IwJuS8HjAE3U0oVVnqyWfruwmbhzJjzLKKYRyURGVwl8BhM2J4lRh
iMQSMvkW7rMwMKzI6iAjB9L3MY1oaBZkqJZCrcgLvt/Po/dUQsZmzS+mHj7Hnv2N8qUjOlMtDHlk
xwl0wYGMR9DzzR6Zw5uHccoo95xXPkIGNPDPfVzifbj0ZJa7ZVz7zpxil4t480S4Ru7NM39250UG
x1GbL3yDeBWt1IeRxa9NQgemrvTQTJsyVLzkFZjh7dTZlu8CSAeqRJxUHoX1eJLoMdY1wJ6c99aU
Vxy1WY9GJsef9tLColpUCZ3R++wsN8D4dZJs/M8QzIDULXTNdEwYjGeyJCfWRu+S8i0ycPoc6oud
secxV7pw33v2iSZp+Y8a3IIbt0ZCeyWl25bbEw0YIYMzXU4Qmv0uAv+5Vv/WCMktzBXgSEliRO6w
Cmpeo+qVCCS+avSsEV9R0SLplbwjzQ7zdRhvqmsCTAq0cc3k0yxcT7a5i2Db+McJOQQ/Dvs6ry4l
M1sZjMv03kp+jwVeQJ3Aji7+haR1q2jXOIpdqvZeEEG4dzOltfQexhp4JrgK/A8TIs6y+qmsjmVQ
85kt5BIT83vIpRkpROSoXvuM40Ql9YKasPTeTW+g0lA1ELshPxXFMpxVgmChm9/9AU+vE24BnKFy
NEffjAJnthDMjc7QC89KUovBCVFrJDAZtDkiKz4VmZU7O9RY2RSRlj5fqw82yZOUVlNSfmaRad7V
PPDz6CWHnPb0pQo2uLpUf0w0g8+lGSHMs7xErWYvCgj7qicOGjhG1lC7oJgwM8V3rVkHaWB2GJYl
2jHuBKDx585tcDO/coyjuwtilCk4n7GrjN8UIz12QH5Ei028sIqgf3snZPso8N4tQXM1XoBvLMhp
CU0e7nc1bQhYMBJuzddnkxq0RV8caeeIqD17cFIRIci/ieemuggoxE4K1FWEQR0fG0Y+1Rb0A9+O
bnV7TJz8D3xMd75LdLxIy2yGtnob67f9J8imq/TBH8lNoZ4NjiH2R5e/sJFdiJHjL2iMuf/6Cmh7
HXv4+yEZbwJ8N3NUlXiRZ7hsjU1TWFPiyTAzlYqrotIoXQrnp1R8LgT006UYWAoLZNVQ9pZj+6Ao
UZMrxWGuYvTvg4pQRniPztvojdWHQygPAE3Tk7wFOWNDR1+TQ8sVY7c8oYWtCKfTQJM+NsVA8Enc
jJrUfIfjxcvZwoGSAKvLxmTt3HSp5Ve0RKzw7iBQKTqMDdSm6lups53a4H+aWiAAyWIu1o0MOO+K
QwB7mJASgJCubXjnsmi6dylGN2WYdXTTSw80mthhwfBi80EdNwCrXEBFFNqTbNqyp1D3vZjYPyE8
ZmNaOB/EV+kO3rXD8M/+2gVKWSoeIPkjbCq+/PPMESCfWDS5Z172w8KUfBpOALkTUU3LfTdmJfDY
I1JJEbzQGHIFLIsxMnknG7DZ9YOpYrs+kPw+sy+XFtVQEy9dfWW1z01vJyAI+G3ik4WfpIXR/OY8
5XXFhAbM6H1+cNfP/t3DB/gOhJB9v5MpldgOUkQufGmuRMHX5IjoqbOX/2pcXjwxHmJy5HQ5ZaX/
Z+vjSAO0mzvkiy+f1zyzsvDvWfEMslsKUBSvOuWE/uVVCKEyD0CyjgxayhrIN/sFXTHLQa7IGZA/
1nFbdBMERmzeJD7ervzYPWLlXY+xNz7ejj12TcZWvgI9meyBlIahhDNV/GFXcnIIbD2sZS26tUQr
Ca1NjEaa900nLGwK8E+cpeXSJ4U9bufBtYrm/MumFpibGmmFzjaMclsq0jZOFCg+XutlzaYclvRE
JTZKe+xXcY2YnVCcthwlOWwmbdD1cX3EgW6bo3ZVMXkEo44eXR39PdbJc67Uv/rH+rsf2dODtWY3
oAoziflc6lJT/AMBZ9iW5k3yW+DUwesCOOemxuWbV6gb7UME8+A+B7lL9ZVndgcm79GMutmasXrW
QaKLS1mU282kJ9kRPMpw+iwXRQnvvrlJ2vuuD/mutXfYaPtUn+UZTagNtk/Z7onZFzZYsmev49Cp
u4zWncQOcSdRonwOFJGY1eTUOKo2oJ2rHjVMg/yx2K3DrvOXmKR24JpPhAVq3HQiBlX8e3qZMDlO
SeTod4yd/RBoG6GVOkiQDHiGJDXSFGRGHfNK2r3Cp58tVTtiK6yktWZk3UHYS/de3QQbyAIzUMw7
XYzdOoji0mzZaLX6hfDjAZJG77NFgCq46tlnJ4E0ZJYlMqB5Sl5b8Db5lX+wBIo6FZRJuWOqpgRx
nSVttObj07Ohrxjw7+enK+POQZma6o4gxTfMU+VfjkHH+wltLD3X7TpqDq5kY3aCOTB0Qiqf7/RJ
k2E/RKreMsGii5nW1aBIH1gy22SZeBNCZLnILVCUs+eQ5Kivg96Y4GnF6mfmRaizUdWCNxYdRrOG
k1mbeHD5fYQB1w8drrrikPtBp8rbnJiYFrU2GZDRysToI6SGpnn4v/keiUSOgeA1W6394a+TdYxw
gnEBsZRI9VBQtAXGraK7Foc1xq4/RKNnGG4HOn877bhBYYBasGFfaHPh10eRz+McdMz4l6Desawl
SlWGHQACoRzcPUijNX9B3LwFjPiuY1BZ8bhT8+G45ARWPIHWY+55xS8D5Ap+z8r3izp/DE2gCvVO
9TrEr1Ake4y5AwffFdkQ68m8ip5jrSLzts4PZzR9U84CfFhBoKHRdaDG9+MGiEa8YZY4DwvounGF
q+SrQnqfUvKyo7SopChtswxY4XVkSonjGUIjvAeR//qOHKPKuZX/Ly0dRMEnsG0TnYrXD+w3gIoX
dQ3YEE/+T8yhADDmmThwgu+TpJvlH5DU3WnoUiK2GRLimFztvovMzmqHCPitnwHk0lOzEJQ8Lnbe
o4vwdRePK0wXxSiEIPVyXSSDKY0nlN9M2vEyfpyw9HBIomho2VMAgDZZlTDpRMBuDiNEcZ1CWEQ/
XgfQaiFfByOO7GPReRi7TYjC+r9wcaEdtFL4jI8SNSWewTAxFMCnUa7OtL2ZKbs0v1UCnC7E55nD
eInlx4QPlIj2yPG/GUNO7H//Iy6NT0qKIwBg9P21/D1h2T767jYsDnWbi00jcux/7Fd/7AMEfDRs
n5yVSnhRpI8EjB035drvVcxIvEwU3a/XnOp+Wz/LYMDN/+ByDIvPq65ulbKoLDvbW4ep4bCoO4WR
ALgrH76uCZFd5uqEBU/40Q41xnvQ+CqTtWxgQF4foqaW4ewSW3ca7MQvE4kZIYconR0eg5ZgK1yu
bEoCzMqzbaXQ+NPd9tLTjX18052TvHcWlgQyzpcq8D6vYt0zkKh74ntvIPSffa88d1QHxbod+bmF
9YjZdyrt089LQYfuCr9ZQtoHubRVU0yqtNLrLaCjAUzGkMrgVDBmi0pi1ejsVoHUgNXc1QIAAi9L
e2WS5Y4UUajY2cbqTmPdkDZbhSCYwqHLlQapnKk4QYg2GP07iNc0zgAbQllgedQIKE8PRY8XnhG7
rYnWaXjrZZFesOolyYmzFEu59W+W3K600VmnwSY8FgBJ2R8O4DMZ7o+bBI5SUZe2YMYO8csPgAM0
zjmhCgTDMkqbPQRpZ5Nn5TZ5lJ0CjoglOOMjoZLNrJAxP/B6UkxbEs8m2QjEUQtFFBhR3BHs7Lom
yGL3u4zynnnHKD0eYzNCYyDdj0zTNyn2uo/FdV+BHBdb380N0ck1+DRQNEWInci+MaejMiov7nAU
YqPxTMZcXfnxGjRNBuaubrjAr5ZHMo5OT9deKWUV+DMoXCsfX64lVZV0vco6meLHSPDzrXwexhNE
wLY2AC9foe8hofn3fVO87ojlu+jWbjSBCIG0jTEkCuCaOq7oP0N+irerMCFF1RMm+3HBpT4htCmG
VI0uxj1wU4jVItEnFH12jImz+VBcTzIa28Yanl/NZ4bZ5fClBwG5CdrUJ2VYEmYs87XarTb46pVH
GY8mgONIRp+W1l0zeKODZrzDo8/KLIgihcrOb4ZFWxwbn+qWG4J0BqF7q5ECqZPbWLmaY1z1d1mV
ij3pM6FwNldFhINFzLuJNxFJYXAT61+arveCqnaNe4T5xpnWv2QPxQoBhT8h89qNZvNtZeNz9yRA
H3togTIefkkIHdP89UpDyHen+H7ZkBhs/LehiSV3wLPLhthdfmIgOgbrDoeq5Zg+ZmUdmYvTQAuh
JH1Q65SE/8eutat6xGwT9aRDtUiDr0AU0enPZlQ6KCi+H6pag/bXm4axDD9ncIo7aWafB+9Z3nr1
w6E48QSdJJceMvalmHHSx8DrsKidYoq15BhbIz9+QIYie0MDd3T1uYSPMEoBcGnlqJop7tH10pZG
or3S3TW4Ai33IkL83GTUkOKeykVFpR4oOnH+pQq3uV8Zae5W87tF558x9QgN8uNbACjR+Pj630AN
Erz9htJk97y9LOoH8fXoZOfhRfbzZYsldpGNr46RtKdP8RWfV5jwAUOqvB8vHoMMG8G5kP4B8ow9
0siEL8hqpvxrEaxeiJmJciMX/6bSAw29AbPr6oKJQ03MZMf9KFEWNI1l1ve4tuPz5ZHg5RN/HxIv
JMzyvHJw+ERngl1Opk8AyQ2sYnnFJGki7oz3WXmW53M6Yui8nSjhlrxUpUKgwD0FwRgiBiydx5Po
NefdC1hw5tgWBgkPXQRtxpHCce5D6fkxBOdCGquO1cRCSAeqDPg/EAyStSs/PIPd0syrIfX9wdYD
J5+xK8ElUMp3CQeeAvSYQpQeJebRzy9Gg0ZbPTlTWcvOBWl5xaQiZ5xhBzRiD3Mkm5UpL4WUnu0i
IB5XfscO6DA9qYb+Fr6X2InT4C/k4ZB7nr+ap9KrVbsmu2nYk6MWSdUERWVhCRgox2M8rVqr6wv9
Ipy19oFngLwHQTtdZTunQI5J2Vmga+XW4D/T5cL4bLuAN2P/JQQvteqAjDVfXnpHex5xPhZrEV/S
zq+JELncwHQW+r/Ii/GDYxHs5k0TmAgYhcLoxGFOsKC0IK6jRFFbhKGFmHKx/xUFaEjkMKAn44hf
T69rRTKOKmn/Il1VMvjyacoF0majSuS0E2ITrIKXLXUrdr6jMsZUFMlR0TKcHoBXNrEdJHgZfB4U
eu26gDRk7OoKzZepzOusD4hJyqK49h+fvT0Ap7GBWvmMMDt+4sD/3TEPdD4j556CFtfwSuCcV6EO
8fpvHae0MJ6FCceZzxMMBNccJztv+TfkBDya3RVXd0kO6xOZdorODBpeeK16aXG8gw1kEGgWc6j0
RYX5kcz4ofPcns8kYTuhjhXIroH3IYDr+5T08pf03P/em+XQscO5DdJDysjEr6syuuuItU7Q4TbA
A4dx+kT79zT+ZVHSlUd/HzrAFN62Tqcff9Q3KPMZhj5xLK46rVjyWiIOggdTwi09SNLzQsF0Gh8k
wvW7Az8fzm7Xz85qWvyZJ7edUArkhJk1dY3AE1OhfIzEQUodcBAAq0j7i8YQqeEcejE48vnpiie+
sC620+H8UBycq9oNWtTyt7Zmc9Ge5bWfRm2OgQ4FnUFUTRxEmab1Jf7AWDH/5RkXoWL9MAC5h3OT
g20EOF9wQloObErep/5NLxp129UR41KrOsm2DiHwNzwkvENRrMkuxdIFVdrJTWnvKMJBxLbLg2D/
FHuwMFoW4JA+Q5bwWwZCwOjHzR8q4cROj1xaLwVjzdjpbW55NQM/iuR2bvbXn/hP/2Q3dOvvfheQ
T7JpUbi97eddEf2tXO4h7Z0AWb/f51dA7qVIgyaRAdTXgo/ASPmi1JWB42ozDxCOBHXrQyjpaP5j
sreA6CKWwYnlu8fn4er2W+3PdROvUOBPbSNdgImcSTrfIdhE7+gG+E0zr58E2RK8TqqEedC77TPW
B4GXrJsbeyFR4efvxaifQYy/Vt7rpFiy3+7LdvEvPb0MrlZydrVO4GX8IXkmQDY/5Mf4TLc9ptNb
Ry4jmzEls96RIfRTXwX0pd6THtORsggtk/LtTFYQ7rteqTrkCpEaAqew1298baDtDzH5KN5kgz5Y
kI5v0pTZJg0o0IYrfTLT1dpvHpW8/g74JcQi5QEEhWfmRP1msFLpRpJxxXHds27SapFCWG+pukHU
/J6q+EkdQBkpN/Ml9dM6XdVw8Ag62SEBF9siD2Kp3kZtdkYLgxMR5ieKJ5/Y+Wqb3KrPxOVyk5mX
60cVgZSMX2aYJJRFW9YkpOI7VZYLLPzAp/8CAKz3DaCcNI6gxs7mNpPSe9xU4LGG+py0M1xon8DN
vcfEWvgdO97CfcUxYThyR2PiKo8icoCgwUhtm6agN97IDpEhWPjC9X+SnAUCZicDZ1VWWGiSJY2U
FopaiUf+LfTSWqDHmfU1d2yL5RHYYdANaCYkt/PT+LcyEGuDpf0/xMexw1bu1GQGKJD48pNAXJoM
WTwBWLZWqxkH1klpsF+5xieHzCecZt0CvBQSobqDLk0GXYo0wxl36KAqeYFOubRgr136x+E65gnK
SMeCrlDCoXRup3K6mPO2yyswg++2BjxJp2xxpGee1e5LWAqH7dGHRPOK8J5mb3HtC0rDR/1xPadI
H7PaRYboioU3P391uTeKAoS/m+IzXiBz0VLKOpFu67xbWkmTV7jxFx5Rbad3c1AQfytFroesFl5J
SnV/osE7EXzmz13hoTav+j0xsXyy1+vaIy9eDZllf9M8leZ7iB76Wt8nrXkZqlYxOZXDN1C4qnil
abh+P4CjTU5sYVtKLoE3UPSLbK5p4AuorM8SYVc/b0pOMQAZUIBwdZBAaOefqxEEofzJ/yXMSuwf
bj4DJIpAbKOtFYj1yJVsaQoTq0SPu70yAOfbAdUPXwbLKPvwWCag1rrnjeDSwv/csOX+Lm+s1x10
U32+J+9xlDwGF+RtDrhJlPvvOEJhOTy/jM5PC+sXyx+7YTOA6aWBxudHm6eJVIe+sZ5gya+5+/qy
fLnBy2GgKVc6O9A7e4AGaD/9aEHSAKWFVfAn21l9/+3QoBJORwjOPc3Hf66eiNRbzHm5eUC39gjR
VXT0jg61WvsFGsptWaV/ALw61ldaZKt/7x8/nZfZwUi7naHduMQkYLLX1eH2eoGM0Xq8BPt+piHn
W+FzWw4FRIM5R2rgsAQheOgy1V3Thxm2LHIoRSTLO4vGBV7QUwRoHnZf1q1bv4Y+upf5plUu3t41
vwBGwQFgVa2k8fQd9eNuQDFmPnzPpV2UxIBPk6y8u6pajPvV3eWmGA5vafgZMHns+NiYbJnbevJf
DQLgxRB4Xk1d3zVZTbTVBEEG0UzpCTL6phuQHmJz34JsSv7lgUQxOi1GQlRtd5bgLngqS4+yQLyT
yzKpeLoUpm1kezKpYvAg8YiNfaB03QWMZEv0LW1KQnuHD19EbkHkQCzhHEBSwr6uim4UWeITZNZf
KDw53GansgdLN5AznyExH6n5typVRffWIQba90p56g8HoWpOosLdIhTxvv8sPcC2UzdDuZAjU5OU
3AjNG27RNz3BHzps6UCiitBN1bI8WQ2lmix1Dm99dnXnZnobnnzltkD9bXJKXnBxcEwgB1UWYP6H
NWQc281eIEdIQtNgV77O+lYR/y0kybv2kJQmuXJ5JSdgNbld8W57U/9Mb3zpr+A7ZNEiWqn4pFNs
LGhXDfQfoA7cxlOaK9p8SqcJ6jMhPD/MZSlhEterM2Z+DrNPDY5ucoGRKONUjPNZaF0FDyeknBGV
1tSbYcJRUrGHB2P8k2cOkm1NkH1l0QbywMgY0UTzgtq9L/wRD6ko/i6Jxmqtaegzz9y4rFb8Pit+
rS9D2Je/Y6u+jtdRjjNRzik7aTU+XqxIfKG1ZWiNHZCWKj0X0bhkqWVLePjOjkE4mFg9MTLBQdaq
pe7q0IC6g+QXxp2U3V7nMjf+9MXx9avqlit8RJ+EuOnh6Z1dpkgOBX3h9sGTQ5OxvUqBy/IiwpmC
iurb2vygGFWttYIEj3jpqIJ9RoWo2ZPDqTwXh5a4g7BMB37sjOrTbmeFij3RrY2MVs1wvDiQaJVt
TFZ2ZMgOqY7TX6Re9hmKK148pHBkrs8AFhdYLF2wHdEbbAJw4Can3gz4tfSglPr2wKnOcVDKEe/r
yRj7KsdxSf3KF/PtZ3z8BT3ahRLgY8AxFeWwRIHmN8ZXzfYAsoWlCk39cxy8yxYeOlwJN/PPxg5L
NzMfM0tEbQEVgbV20DMqtUW36MXeT8/kkc+4yUkI70vyYvtHuMFX4WzUVMWSO/M05IhB2Ak+GErq
ssN6ghPrTrAOAD0kx9mKWg+TTGt6LAEX47xOtdCO4OGFQ56UgQT4j3MWL9koZLW7kOg7zkaHcdEK
PRvvTnvxJUTiArHX54d8hDyKLYU101zlVtOO9gvuts0WIbR0onn5VWofmwvcvm3Y6V3qnIYW7qI2
8fmd9INcMxNQ9dmDcwprgcig2FqvCpfNKtvPQgHvmgn7ene2cXjqSnklP66ay4KnAFu8FbKg57NW
BMajdlLEp9iriAiqqgWKubhw4N554M4MCtMJod1r92rlvtU9O2sX8Ul1D5NFw5Klvf4RlUoYK9oU
EnlAA3eLXRbTDbDebsjNjGJ0xex+sIZ/OU6ocpUHHiBBX5Ml7j/svnBSZ3b2qKhcJMRbsym20L6d
pJ7QiucJpyz8B+udbK3ZR8p9xWI9NhY4dAr1ZqzOZKck/u02rScpL0DpA4Gjj2mKYf2KLFTTH7cZ
ja1+vye28suMdks9tiogg5KlO+bi1WmgDwC5DeOzoQCb1M6K2WOQNQVRRu3xoerOyjpIKx+yWz93
u1424H0eZdHJTKqaN0viDRpyLrbfJQVm4/bURETS7g1sW68ws8bcV0t9/H778Rs/N9f/xkv6dpQr
04HsSaUrOwllAhXTEG5R8ylJZRoHX/NBDMcq3KpFIMmbclwZcwkORy/mOgjCA6zza37anQUL7olu
bhM+waokW+j/HZj07AwnLMeNeTcmdq4wP6sPZmxpm+umjG5cE2DaDKAUHryOzyWGXKI+bX0KHXiL
ptGcRak5MHD35H4YoiR5V3LFqFqSdYkpCr0/qYAgQt9R8FLRDvpBSb8OG87Vdnu8z4o+k8LIwfvD
eFkQX+pbE+MRGUCXysq5rVW7KbWdjiqw4lncyyWHOzTJ1cHsu30wbHWUfKkDTtVVOOu4eQn8inEC
mvY2kGT2T1qqDrPLkRK7Sum92tj1A3JcWpuGoE6K4WwmdUyU/bgsp6EZ0kGFWlBNrI3UgHiLwm3Y
N2dBE+co63oBYMHsHEbZSWySBGYod1mXBI9jhsx1C3BpWmaPWbqQmi8V2yea5rcH7Ds0sAu/NZux
frTH6QnGdxFaEpa5Q1w6nDi2qj255ISugGxbIc1SQV0NqWC8yYXWeHdvbCpYslCO4Rm3UgDYa3+y
dqYNeEyIVgrgJuwp9PrY8rYNWDvxeDW8MDUt8hGdt67CAxk8NoZty97oZV1m9ByRRB5OzJQCJXu1
klCUZcjxLPEipUuZU9QnGCDJYC9UZeNOljZDVp1NHWvziC9f6oYrlrJyJRKuU3qYKPMVWtmTjC8T
2BD+ePbap2PZFeakANw0XiXMeg1HjMeyuOr8myDo8mBqLxBG4fbMCwGF7hZ9X/6a8EPeSeFpcLCN
HEZZaS/Q5+m9OehIvx/u0bCYskUR6D+W9FOwtEjm9zmNBI3UmYwF2n37OeAm0DMSlQStWU/8+DQ5
YyZJ5NQFsktiQJo+qOQJJf4BzpecTNXfF0B0QbdDwz/SpaCh8QRyZlq5JoRSfluIKDPJKLh8iugr
MOYWl3oX2oR1pYDatQfGfOcY2lHGZhXU8apA+8z8KWtPVKC4z1A7ZOPqh5z1wAsDyfP+oERzq31p
nvoBe1hCH+feqiRdKuT5/T3nu5gFfuMd0Ekraz7iXhHJK4VItbOGhWmbZwklGkV5z1Z1nnn5Yop4
OvFOV9t4Tw60tG9N5XqYnbuuqTi6Kn5WkW/xG1PKfAb6zcbon9wCCe9b8DmMIy6GQBJ4L40TbBMf
hObVFkl+cjUB3po675CyiB2BgkWQNX8rVx31Np/AecOhZ1usvGqxLdvHfMQhS2SwNKhdLAZIECz5
ygwUiH9ZJmBCxxhvzzCX9uhXkvbUK3IzZ9LAzDYNxBNsoQhsUhJAXi2BqHL4+43zFtuw0ybFIRhz
ezunrrhKZU7kWunNvkDxPPgMf5HjqGbaMAx/fA9S7zjpmXb1dKoEXbrWvathXY0F4KcoZHB58V1G
OhzceA07Y+KL5wszl/6bTXS3Y0qbeNaCi2jWLQCkRx2MEXjkt0bgz4CgIaQ5V51e7eyNHOt797hS
vIIZHQoKB0zhxpOgDoPu+33bFkphgzqpd835/VIcHDdqcJJZcd6A5Aup9Og3arf9blR/1LZnlyCV
dccjLl/TAb+5VI1YXup8EQ90O0TsW6WnseeoOY1PDEclrvGm6TkmhYdb5nDZ5lQAiBBUs6kvV2D0
IfRNaCX1iEYrbJk9ftwFaCUwC1+qgBW1k7qoY2pGWFW7jNd/cH2Vw0xGoDqeRPukkXbKNBf3eYGy
kz+9E+HH8Flwt7IoXsLSci/AL5Mftd6ELvlpmPnWclWKWdb+zR8+YBho+hGT252bOfZdQqJ7dHIu
jqZAZtlSXJVNM2AlYfZQNsCOQB7nBCGXGF8yIE/80EJ+VDKZK1MtlLh57Z3mIa4u/jqssAdX6i54
yZxFNfJRTRdGINmp+AaRc8phs8dAeYmtEOSG8tyTb2Ppnfeeer1EGq6CWsgVi1NoeHtxPg7t8pdP
aPDdIjTbOtVXmZNrlm17NbxLXZ3uQK9E/fL2W6EihbmdMUj7Y3km19FgKAHTyy1ApfGa/gRTCB6q
895X0Ecepc4QKymBlx8TSdzWft7yjxSczEv19F+q2I18/v/YOwkCS1Z01LH2e8FzQgvw+aztOKj1
dO+0l+6OuTZ65Zgz1aYZnl0W3bYaAvwnMYBHKx0K2FRIat3HNbVC9dfgBKl4kMCu00ackQtpBzUz
iINFp1H4KJZsFHAaxIugc8dPOnI8bVPBexTesieMMFmHFC8OyEq2TW48GnPxE0k+41u24CW3ulsm
YgsMEvPWsQb5qITUsqvaRYPWoqt+CM87pyqZgNNL9ZFB/v8HK5PbbbBe6zZais+5bhN5SD7wHqj5
7mjxxfABcl/3AO05Tbqt/UZHFV8w6qnTCTUzUfeNymd9DUPY2Ycs5VA2uLkLsWvgrNY6YUe+ndKe
/O0diPx5H5Cjj7az3eBA3XzhfwLjVrJr7MHzYS3uTsvnh2eK3FlaThdazBwdTKoaeiOl+UtVRdau
OOryWAOib2UcnUzhexqyI67ZG0NNar9wz7cL0R9i4cQXYXhv8Yr5wzZKFduMY6qhU3+sM8YuleUS
z+SvCsX+ONWiiCn/VCdEJfQJdyN+ihUs0z+/6x1FpMQLKT67/VN1lhh3+bNUN9pA5Ge2B2Ag6uRY
YWAF1wMKcXv5bKncBk2S5xjDNM4FH4ffuxatxVAtF0C98ecV/yT8UXQOMSlqsOfRaJJGoH9YH281
G8pK8hQ82GEh2rdELF7BRmfvNt2E/y/yqm42TlWqoYKoil6kRAuiiFdjBgfTrEaT6AzCoM4y8MCm
qrSOGft6PojMmAQz4jB5uZx0bjje8QGuabWZWMRhF28Q6O1md5oNhPeAzi6edp6OBh9g6gZbXvfA
VJuEXWNNy8WzPxXkBWwBGAAHJQ7Wx7MiDN6yrK227vp+ezCI1KW8V7KNyCSYG/GzYi9xI1/pHGV5
VPGkH+jQkAuEI7KcBnqUd9uSw2ObN2g+DVXfXa8FPpigIvwDVEs6qhy1vNSn0HUpQ9O1+ccdVB3s
UBBCsNqOWuGalIaWz+I4lBWa2kbs/JTMmUb2hFVhJERR/dp5BB1MGp3t8w8muSnrxgjwAh6jV3/9
u6gGQOp+skfWLDYNgW3Vfok/nXHxKtKenOlKlYUHTsR7cbDc5PNAUEXP61pmW58QmQ3IR11KnmxQ
FY8prbZ7C4oQAfYHba3tFDYXuKS+sO4ZhYUYTLFTFXRTDa2HFqNekihG2oVoyfd1y64VQyXD5sUe
Agz5AOCAK74l/Yvw/PhWVAJSHViVfasmY1gzTSg9uktQjPW3/sGzs2lpremhpkE8IXZbJ/Lt670A
4+DnHwk+1ip//TwdsWw45i9DbcUHmbhbboNwUtUH+3mJSf5F8ZQG0oBG3K4aEIXiIU+sJ6cessrZ
hl4n/w1iEAYMp7Y+Q13W9PDw/HgxPUxdg9LHE3uJ9J56zITjH/zVojvd+gaMzdmaJc3oXSUHy0o7
+ouRPt2eTT42OA/HsDMiLpLIIB8S04sRa2ypJkYWfhzFFo86r2vigPXrfDXUerlXGg4reQQp8XCB
CH7omY/DrtFdBiZCIe5KUKoIfYD60o6/u2HILORHkHgzUGmGNe4F7VXVinyayZJqgnIqbySEysQV
B1GGQV2JrItzR5cziT0el4mx/ZHAzaEbd8NHdA0pYoqOCZL5Xya9MKVqnNxPjmqisQR3cIQb1G5c
qt32MUQ+W5OdvhVxs+JbPmftoQ6qJLfhBGiPsHiy0i51BqV6jJTd4SbHBHCbdAEncpiQ8Rcl7fYa
OCVNXRBQ1ZsMxw+NRvG3z8KccAj1ANms9RvIdjmCTB5S3d0WZW5Kh98ua7b/0AbGkHx75Es6mh39
0nWJlK6QnyB8eN3VZJJDjvz3dXwmpE8JRNNGe5cC2FZrnUqKMApM9hljXRbyAl/XNPjNcBqN5qcY
i3NDx87mnqxWvly4YhVJeMj0WqduT6ukGgECqxZ85Ha1pmw/qdPaGHj4OGR4Qgz3bgt+OANmnTsu
kbePKSdv2pX3piskUpkLsnUsJiGW5TPPUYtw4WIKu+f2rx+B1gta4CjXNkX/S6Iq/+ES10eOvKP6
6Y+rKZV6+zbAa7qvBNEgg1sMOafOq9Yruf6iSFjxYN5cyKF6ecN1atInj+yziAX70Ad5YeHRuwE1
tPBK2D4l2ATZpB3wr2jCX2iUMXAZ3F89JeP7vIvOkecqOjx8MmL+30v9iYpuYwqbrITmyNeAEpfV
Gus1hb3kXagMDd1oPPfRRttK34u0HxE4Sn0CPvMv1bPpLUxLxCJbLVRd1blwfUNVwJXlWcBLktFn
09QUujmYRat/zQzp177JBv/cPfe5EEPcu8Nl+gtshTW17IEpROHE65wfqAn8NLW6K9jMiLZAHAVJ
StwnlCDXLWwFyJWAjAuhl9RosO1ph43Ay8lLpSPAC5CTV/cU4j57Vwel2iPiDNuFhVDGhV0aXFYA
hZaEFVZr5czz2lPEF3Injsj5LzycL0aihUNiAtD8Y/l0JnVw5GEhqcZTL9QORILz7oJ82rW9j5M/
da8R0o9SBFv18uJLtcslQ4/PGHvxIwY/Ts/iY5BlK/OiigHGMAOIhKzZqKclyQ3UE/4/g8Dy/Uci
X6lClXRp0Tf4oYfqh6ckjKMdkCzkDnws6UcXs/cJ5y6T/Y9HaWRNmimD1ZotqpuJ0L3mdHcEuFWF
jfb2Uqn90uuNzGvAyC7FZLXjgEnVnEWm4nEQRlZBRjbgIMUVnrnNtno440L3ClKE/dswftTSMCAd
iVW2O5+/TX4qMOHxhB+RjakdI3PgYRD2ugRm3wBdhZQB8WE4ofzIRodGIK9n+yFmOv8bSNhrPfzf
0WjunEXElHJR8eDtzR1BaVPGThYOxqQ6NcYzCB6nsbyuuDZcshw5HWP4Izn4ZDbg/nt1IfxLHqsT
gY0fkbZeNyMeZsQHMKPTAOQxC3Z4MwXd+bIWfpthH62KexXQu1tidZ1il+UhzM/wwwA7jQC1IltS
/4vg+ChvTv66otPT3kYX9p6HyzKxjMWDdhyF32TOMFg5GJRWvBTYmKnnrhszRn3IrlW78bueI1Hv
irstDji1GpRLIHkiGJv3R5aX37u3XKzgTaNbWPsnKtvI0EHpYw6uw7B2rAgOtlxt22+M+IO/pSBb
KeQcuYuU2UUZUp7A1MiMOlV352Zkn01HjRl+lLwr+Tr0WrSnPVgiA7WM37xIuR6XvFn8cKMAYI/q
21cgZRdZ0Vq/aihXQ+s3ILOrZPSbm9XfXPVYz4Uy463xjzpT4GohbPgf8soYFs86C8d5i7St3PQj
RI+3Jn4Jv7Fr3BgX1S0d7JMfSjDCfD2Acrg7up3ta223SN/SRznDinpJCOYZO+oshwS0T3GMCite
1gIQVBDGFf1TEVoz+Rer5onHFEmaHuflgT+ZkWpFmXO6P/rjbVEQfRCZ3kwIzzLdw9ondo6drbrR
+kPN8HJRsIlGYqsXhW6frQZr0eq/sve7qye71VjOKgYQyvvnqKC9TzK52Z1UpFkelOKq77fhvH12
fnq++J4rOXXrA1Ow6qM3oCaPMk+f0iI7OA8vG5sn3RgE+gstngTB+JloNVX/V6C/Xdlhro7ZWf5/
dio9QEJT61OcooZrQ3BdomMfOT1y3Q3pbFOKceJQQrSRZI2FI3NY2Z5smDDg42lbgcF41X0dcBWC
1ep/DEC0D4cMswvemqrhk34waDdfOwUVhwPqd1AbnR6/kItWggl9Zmi2xG1E8IcRLT01chZuu9TQ
/08Fr2I/6CdkaYnp2Erx8iOmEZ8XcW3bK4SZtmmL5fQYbX5B3o2wQSaDcQ5mXeoYoLYgHx6kf+8X
N71NLsmN1ZSQOkO4INPrmThU2jRFH9yAPIFP+YHJ99isIrMmpCA2wO7NN0qE7MoFyD1qrSak0OUU
NVg04aLZwuY9jTMdv8x3va52sVzyeFxGlu+dp97oL8EVxEl5hKjgA060SMUOCQeo086iOBLW3cg/
MIxwHCrxvHnhFBvEmstZika9u6KbMdl2NryJPuzTFpnvWTPaSteOFj93ky6pI0OxjHrTXewgZ4NT
RUnGoSZreB9aWMd1w7brTCFgunIrYaROYom6YZEt3C5lzRqMS8a37iyhJVSZjrHkXwlosNes7w+5
icafJ1vea0O2/VP3/S7kkekQdLLCKLq27dLD9pm68IXhie2KHx87XRUr8DMadealKXNmWjSkkZPJ
I6JBM8yhIv7CAhQvrSteQySga4PGMryGI0hOfgZujZgkqKt9z5JAIguudhmXggdjqBA2OIrrtdkF
E4eqSugmembWhqdAcf6aM23Xtjh/Wjx7Yb4avwh+ux75CJISkJOysLFUCsb3/XN9tMM4LjQAYc2N
6jB/a1C/7y+52uEUvjpcMFKzaHulxC3Sd/++h9+iZ/q6ajWj6Dvz3PtE5c9LiPvDp5Ybmg4Lv7Ap
VczIzFl8dgGIMWG6FqdMkArgh7u4sXO50m2bmY3Ypv7aeNaRyGKqffT3CAPttkQuJTLZUXZ2Bxvv
n6WES4r+iGLlHRjf/TvihmOs4goiTIINZ+3NEstmRHtkGQ7MaJGhk8nvC4yGkr5bJh0M0CsqTBWd
/oVxo8EmN7zq65a1SuyAh+Gvju5LoKpuxKMkBORU1E+k90/cfCjevkj19ScFuVkAM7pip+73MaHd
C/0BSdVb6udJKq3UvGJ3uHHudK9EaEtypFXhcbq22H4yqoGHj1ka0hlw+E03wRCL32MvCfnQhkNx
C+N2NdF8mMK6UCRHz7365WLU0IZ76kM8XXWJvMh4j8PZDZtN6WGkz0nXTNMOChM2yb/7W0tE5YXU
n90X9hfBI951ROitrExchuHB17BdE7aE+S0k6LPrlWw1BgDXaCMhykg+REY7w4jEqJu/BkIhxCDB
SnizAxhvVOFL86neYb6ZKO+KtBSgkrqYDWWSlN/K+EuuP8KKaNBisdI/wMXe0sbWGi2LRFRVzHd1
77Y7uxVnCD/OuiRj5GYvPnXURURIuz5/hA1O0dy2+iATqRCpji28el36eH/QSN+yQk4i0CCf2+WM
uRaQk80DC1gLhYFEdhMd3x4qOMY5NxcLG/EUMqrOszQifOcPBExwOYsNh7oocjyu9M7VG8WQ54rT
dji7lWfyKHyPAlxwqQMquoQnZvQ9/ECg2ZJAfV8uX5dkoz+MVp4KfJJnRs6EbYDZZNV9G5Rkz6uT
cma8A32i7bHkUgKdNeOsTjKaUp7AeeYvZNKvoOfTtRTXgPggHQODT3nJ4W8wkxg0QAgI7t5emsVG
IeeCQf2AVceC5eQuB7KHn8C7tJdZdCZNisPZDqwLzTstyNDxdIr3QTV73Xl8D02yNKGxl+/btLBE
CqDUGbTrJe5NK7yqtp06Uxp6GcSpo7hn2WVvRLNfgz56+YTa0b4jV1Vw1RGiMEdkcm4w+o7kHk3m
wiX9eGBFE3ai5lcCkW3w/QJJvuoFCrGM8pYz2xLcsE+Sg7aOpN1pukjA7KsgFfasS9yhFOBkC7YO
y3VimVge2nfYkhm2mmijknyCPHV2PdQkZCEJP5JnrESKKtX+V3cwd+4F12jDod5t7Lwa9ikap3xw
nHPRdRzYtcKUaZu51adsrlfbpJjW9SOl3FHu4WIbI0cOvTElmgxL6R59mcUEiuPWqv/f27fZv2Bv
NSMMdjLjOrXfLdUtaRoAwttU0PO0oWPX86KRphFznMwrsdrCnsm2ywlJ0Ruxp6MmwasMOrIUHnBN
yxbA2uKYZO7DRktbeOSLpAxnEhRiKmZZKFZlyoPI3EOZJuSU5m3z+76hkec3G2AiZmiYZ04QChO+
JhaIzpG0P0/sCHiie83g6jA96z2n9I4aidk6dd5cOP5E8jC5HeJBIR6m9Etk1wxwBXWpMkNxj08x
GL6kNYyjByEyVTI+5IOHQq8vUDIAhusd+t4uvZ/zNxj2+kqqStyN3gcjLaCEfrT3h8bGiIac61TA
uK2oSoPMTl/++aa5ooadSkVWu5PlC1XBx5Qv31v9BfBKDzzVficqtlSQP08Oh6T6k9fVOlZhTub+
Z9M8asAjabDS+ghfWqfE00J4Vs1U7qipC6IRfr8etHbRYRHnv/Q7f+T6p6MZZkYlA4Bj03K9QxUM
odTlc6JYqPwj44wyXbcWpKSWINxnIIeNT4DXTOfbCaXMylJl5oEnlpQBSHccdiLOCDBIcD27teah
IYZk0rkrnhngDaYS4pslBMaheATYEmGixgrtFbMfHz37opA0nlXcA5eQ6XcuXOVAFZdwrwTCOEJf
mubtPy0uKTMhO45gM4pB/NPgxdh1CjeOsC+ynReN2hAxwIfe9j3iZSRm7nleTxzcccOVcMOyqwiD
v77OkyzxVsIZvriHzBQVFwzaR6NiFd9xL0qmyjF/73UROoSetuUQ4zT4eUuBYjlBWnkwYRykadNz
grmZPS0qXRPOa8k8ysoubN0rXyxzcM5hUaez/pQgbVxz40CXrF3/T32/wvwH/nUVk5p+zPE3rETt
eBDSWGVoxAQtwwl78GmJ4hLSreZT/3ILycQ5m+X3MY94/K0UuyOegSOSiI10ce28H5Ed9xGQgt9U
A7IpPUqm/0oeVmq88prHoobRCI6M7MUEH/Y+uNLMhsrjS1UMyTZ6OgauOyxRYzv64bf/i85T9raG
zrr5M62LOQ6sfplkudg0VkdssiQuNSZ48bJoZ7/7mNiBI01ogp9qDFHMwCpzR3JQoepN2Xn77ryA
7wiB9qy+K/02MxUKcKEf6w6E/UtVqCRtthfUlVvu4fpZrjM+zf3qsOobzi5lKr0Bzv0qSqqQDZ7V
HFry46Iw4tkImtnJJ647v2Fn9IhYx+6WcpOcjZkUXH8FdGqcAtsmlOXFVIJ7miRSMk+c/8v/w1GY
WA85cXelkvTdTCgouX7T40iN+eEN3zze1JdpiTCdmhngCqtJf4hYF1QrAcRHvI1Z6JajM1qJZ8LS
gvYpaXRxot5C8J1J4pURtrE9jjnXqKgAGsomI497h1nr1c7oLN1FShTlvQ6y51e3B9WwE5Pmy3h1
1haQ2byC9220uIV5tXmWr0oZpzXktpf42yr97qKoae8neJII9XQPOP56VftBtDp1fvzP+OixF/BE
uYFCpU1CV/kitivJJgxulMmBtwbdU6AJVmvX/VMqrP/g7sATTIrfvsJOlZcT+6zQl9NpnggjXt0U
+s7JyeavNn7mYEfopmwsAmqJO1e6cealJ4LNx9N9JMFh1ILH3ryXKUHNa5DkqQSUMgotZwtowQjq
fjGAEgIUL2HG8ZHawnUGfPLXCargLY0S9zW26zVXF77f5TmWTqVp+HO/eNTD0K3AYmFcwtreROpY
oYq7u2pgVmtQyFYwqWfPsM8n/rmiqAb3t79+Lcq2OPZHSM0T4bPqOp3LrHeKpVsSFm+WteFOVMso
XXyvoH5BHVuZoO6v9FPGi0vj9VkcXtT1gBUCa0DRYCSgpvQEBCKb+M+UCwvRKcOU5/Q1M+leuL1t
5IgANqGRz6Cee2JwNrsKqpHbSnuV/68F/uronSwkv6EWKGd8Nby/QX3brtfCUhvdNOkfZ6kywh/q
+RnCvrLvzuzG5aqghyMI+lg/9dZIyBiCmc4nu5PcL57w1cOnoi56xbRw+fk1JL7ner2aQDjS1tRj
RLHl2Qh0BAGfAQJUEPIYW0JA0tOVVxpXSMPve4B8rd+TvbtAs5WOkhMi5Q4gAQadI9Q9INUVLEhA
sPNHjc2sdQiCtBzcGyxsPC3hIpQUoNHoJbpWC6sudjbmBqT3gnpqmMg0SqqyjqgoBOinrioPgFdu
1pNXG5Imv7tyklqS03FY6/084005xonDeMzx8Pfaj+1XP9tHcx8nuLbwRg/YFU50+5vBf7mTL0x2
2B4ppluGmSxNPMQjCyOMJPTSQ31S6vof4apHhOe9/DBRdWHkYKPa5VMMvx1HOBis3NP4eR7+ym6C
EeODjQ1TBmI/djJxgL6m+kQ2l/1mqTTWovnwVgWflPkA/Uv463ufJFXfRPOoGlak03wkqehdEf30
ot0x0yFbKnxq7OP2714kOvPb0XDoIQAVmNzaUoi0wSJ0qcQRuaJdcY1qcQfKmZGPuXeZdL46ULmV
vW17E3MG/bCJacgs50LbQuG6Tneac9h/qB1LdcA5vEErvkCWKKX/RluRTc8bBJqhrXcQ8QjGszb6
YOxdW6HRBQjoCMJjK1UZTJTWf/QvJ0zO4cuwr/zFY9vcOhBFGBs3nW1l+fRkcXlGLUUboa+p3hjw
gB0A8YqHt3mT48B6wWzpd7q0y2IJ6jG3OM5UnUyKWG2bLByRkolUgARCLRAmBCO382JpYnoLsngQ
Olw6u5BKlnjFh6C8PRtLPypGBkMn2rcL0ohF0X2YcdWxFLWbMNidGoML+WFga31p+4dMzpTQdrgx
ULb4bHMouK0wV56VHy+v4m2/bmsKHoBOaHRrNc7xgItviH9i6B4wmYJsj1kdNuOC6N2p2iuegU/T
Dg6IStEp7DHJxxPP+G2R7cxVWa67kQH6LljwcuTgH+wE5NV899ys48APFPDEFQQ6GbBp1h0mUlW/
JFsY+ShFAHszTQj8+5nt45TfoKXCX8nw/9c/5j4VT+owlIe4yfp48Y4Zqwa2zP/PXWw9u3ZzmAqa
nTxhxyJ2aeyw+oGTzCfAfV0SUs0akRMsBIkCgk4jNIPsNK4DUbyae4VoaI3JwkbJ/RDvuPUpnMf0
EE0PZoQAFdvutZi1uaQeYpb7q7EG8hm3dh2bZmblVXG22A5iPDMD9y3ocBMhM1LkdR2OdYjL0R6Q
4npfK0HG66m/uAnFmXv9kvYtT+jBPEWWjvopzskqyrJs9So+18zbn+rN/gjxAdNhg+D85GcPnsn1
SzSMvqwjDcmev7HGFz+DSCETlR8poKVJzk9/+qYr1f9kuUKJyqc+g4r7D1paHuaHLEOc9TNW/M73
2jF0enWhaQMVqiggpRO837WkORmweDO3rf7c9BufK0ttyVjuE5r13yHn/KQ1tRlGH2yAv53WEZiX
oVHZ+WLb/17Deg92Xv3qTcVKh/6I57ymAI+jkjwX/6lkx8OuSgUxUMMem87n5csIgKx3fUT9r0Ya
+wtH8JUofHYN9v18OL7Wvj0v+kcJAYO31y96CSN3CH9fhSoV2GuAzRGXD4doZsNxKsgHa+5UIZmS
Lg9lsSlAWFRhEhHqd33aQRGR5tYXIL4YQN3qb5mQMeuoRSBZcUP09rtLeAkta6qykWZ7KmTg+I4D
jhHwomwXhfl3hgP+FfRS9KIBuL0mQAgAPCaDVk8fQaWpwKMyze+pPDCA+tJ/33P3c/psMGdwOjMM
IJqfM4WO3ScFAVv8gr2T8tQZJbC5MOcBHS4uoLLxb4/eOaWbLJ2xSBQ9M83B3wU+nxiqsbDijwlV
c14Xe/y5P2RGNbGxyW/OlzhmZAjYU0cVEbGMeJ+vPHZC+f+MhNgiWAIQnk6m6VfNXSO2nhyct/Xl
Shmp3ZMe3LTupNXgbFJrq+Qqnfwx1SUzhGWjuC5gSGzho3ZzLl5gkTEP5KBZN1L1RIaeqnvsBzZW
AqSxU5E9xjuOrYAO40KQveX+HcX0e0jG+GCO+mzn7t9gm1DwotjlAnjcXoMstA6JjLvnHsi/PzPx
SP70W6WmfNGzLx7YagYaVXhgo36kqOTQbB/45DVt2DltqJhWDHL3epUsm2srqgjF18bq1VRONLJ/
UiJdVduW0jaQW/O3gDtvO3ziYVZblBCCsTYgP1o0kFBH/M0XbGKkjVfeMDXJg6shH30CslHhQnPo
SMwLzirrOowtgJ/4dmJjeUK1SvcpQS+h0zVAUnoxMb0nkh5YJHEWajf81bE1t8QhNbM9kU3JvPpZ
UvAgSlOwBMwZ/cQFWWRmChJ4B74NGKT4rrfYLv229FvilVJWVo22NA91HAMPWtYqj2VGdqsrvFh6
FDg5XcUrHnPItMt2+nXx+IKT96/govfZbyR3M2On6HagObDG9JBYXBqbJFdc2Rv2FQWw8xxiGvpO
8qD+caM5KdbgEj/cX22EIfxgCq6gRKoxLDjbjdLplZhFch37s23U9Wm4Yb/jZ02jGXDRBw6cyte4
B4Rp1HoPaWxcF1GqPex7Uy2KqyKvgS5LgrrpGc2lxrbrPSA8wFCGN809QHmFmM/fbrrHnPN9S69l
7l07eJIWfz6KZ4hEe/JuoH47Gasps6KfRJ0WoqLPqimW7FZby7/vql4VHY6CxeJ1yc7Y48osalhO
5yO6pxhaL1ZLuklJkzEl1szL/mhwM1nD67/kths/PeToXVNr81cugTyq5kXDmHe1xCcthrv0ouiI
j9awA3MYG7PuHRQcStzx6yVCmweZ/LcUwp7Csp/gg/3gjx10E87KKLW8PITmVpeuMB2e9nQhHQlC
c5fzY4+QfAAQxtUyZUUVTi7cGWto2+UWVj6SrT6Xi5NLuX/6L/XWSnR4bv2IPc1X2vT0lgabEuAY
b+KXJEy2MfUCx+Fekr4eN3ODTWK+/W5EgEHMLNV4cOg0I1LeUiiTeR5grmijh96to9ROtK9UJMb9
J1Z/tYdDcvf81U1jOmkiTOi93Y7MqLYc1U+4w9k8ODDPc4I3HfSC69FBtV6C6w2Qf+mVso/j0JlA
m/fHopvP9ZW2ZIZezz+soKuDqLfZTebfzzhX7wb3+8SDu67a2FDLeml19W8Dcx5tZ6f5hO797vXy
rEGa8qyK6GWXfK6ZuXC7+WWPcnl9sbgDwzyR/1VU1A7CnFyDCZCdIFjj66mqlMt5UZm/I89hYt18
KwD2Fu3OzVHhk6Ma/XrwwOv3UbUy6bWO3v25A5e8Aac3Jt1L1zBr32D3wJ39fIAL7FhWXFuKTFAw
v0dw1Ml7yllfXws9pkdAInQtuLOGs18sFgaKIPVt/IkQq+w/eoIKj8A2vtnt/piyTQSLJG0CQbjM
JVmE/eqNabqVNdEGlqK29tgid1JqRjrUtp72QkOEmbjOYY8kQRplTt74l0SOiA2V7CDwkjFebHq2
rseWzk2S2G/E2JhOb5FkRe2JvaJBYGFSNBtet1YP5Lx2Ixnd3jTGkWs5Q9mDGhMG8dpSbXDPBka8
rzizL/Mew8omn258ue1Mc49a1Kdl4dzyT1DvR+eWu4vBMW9D8hZjg3RQQTdT6RN3IpuUwB9vX0tc
XEmu6rW+p4sFAkmGwbQIpl0aPZnao0REQmwAe3eDST198KQ8y++AY0qF3oaup5NL+lrmC2avxGIW
/lcWBAJTxfHeWK6gJ6qGhgmjndTu4LgDx9QYTrk/67+a4eb14X+60UWI4tOYxNmayV7NESNGp/44
soWwbAETiI0FIzDtolzSivEIpmVW8m+hbWWiLEOY8dgJVTLOmKCvI9G2AkdDKmMDjyZtuFPiwF+Q
o6X4oLvLr0XJPPSLV0oRbvF02AIsRdZTM5wSuK6QoKKcJRGPO5V/7DLYeD4NCQE2nCRUDkTO9Jqv
6OGhjsXgrd33/fUe13j35LeyUPe9o2o/iD2OlCyqtNuf1ALKNVQW39I4RqxD97JGEykpT5to4KNz
G9bCd4uEaeEEOQGfdjagbwOJHDk2h8J0juuhaUYwlTi1WfN3xM//Tdj0T4Wcgul14iJZKMHATERf
RjuyQBWOD6FeANPTUH0FQ8lFudExJlwWDORVcfGCACwJSE4xkiJSR/MREFgEgvVA9oQYbCiRYMRz
FK39D9ofKQ3NWpYwSV5dWeUZZhgLcmJa6mryYF6d71YN5DAhdrq22lLDUFjE/JAQCTRg21QBw2Yl
BvYqaVvCKwMUYVW9Z0R9mAmO/v+QXZ8fQDcwHctD+ZEMR2DUZQwgAFN4YiMtqU9N6b6ndwloqLkw
MqeDF6SG0QpLNmRF0GtgGm6Ou+qqXFTNKx0iy9XfDAtzHR0ySsl1chtiWhMYiA0zW6nRcqoKhkdn
IxJqb2r2F47LSWxT0E8okSb/KHjhI/nnVg37T9irt5AW78Ex0zYzrqa1mUOCwr2J8JbokQKvDkA7
LTC53rKT1KI6RjRPZz6sfQBxX9wNJjDrH4BBkSFL3+34c+zfK/pMMvxCxInlEjkl8wIF7vUCjlci
bz0IvWtjwVdY4X1PFrYq6gEI6jrfET2iJnQ8p6bpgJ3EtOaqCEIL45fVAWNGbif62MC4gEZ6CTQf
DkYo9MElvKeJoX72NmRd5rmLLyimue170wjiclIgDcudR/CyuTvugfG4aRaMo2lCnNM1cMOX+VKh
dox5SbTPKXJ20br0ahwiAUTtkcY7RzwNbJVH/Mzvpa19WF+M/D/QLLjsYEWL/JSeNgnKt5hIbug+
HRWbhxxVK6zGo/foih2gPzG5wrrrGhSh1Wa9t0qHgjG2E1ZQVZLTb1lSyRWQgJespYH5G7l2Sz5M
xy0WKwRKY1qPmFK+CnjsF3koBWWwPOljDMHrN3cfcLyCqYmAAc+F1PjaMtPwBYLYB5ZFU1LyeDs2
nhtnxNsRFXvUSwW0lnCIZYSVfw+IipJtcY9wpWpiQ9Ac1ktoAGOk0yIkinH6TJ57TGerzcvtworl
BKi8rbpuH747YwyKL/q00NZo3FG0Gkt/T5bpTg8tW78ES1BFTaf1TeV4TADdXAkUCm1zoE0IEOFz
MqKhd1h4GlGcuZIxtEAG0ROh2vdJZp2UxrNy1t9vXViXjhheD0ZX9u8eJtiVI8ENqaf7+Oe4/7Xu
zIo4HSHIWaGmcuFD5TkdK2CoERL68+J39RZktywY+NSpEl5oPWBERI/S9nTWkv+s+rTFtGSkZwkE
18fEQXox5FsU80Ie6hC6ItZoAvpwylBnBjwDntQxTtPBhK1LrQF3mlpUV4xRCRLlpKhYF4qBiXRu
uWW/NuCTQq5P754XMyxAcy1ves4FTk/tDVB+ZbzIKRX9OeH2MLfHMhWTUwr7+Hi3wOrThUpFSepi
LNIC1IZvKGS/ELO0dT4fiUtuVFpWOABKUc0AMeRnJbzAmJ2aYTM0SjK6fPyyD0+iy/3/Iuo65rO+
B/2f6XTQ2/ksbxy9uaRNglCvfuc4cGbthneJWZgL9K5m7JCGMbs5lFT5rITg+c3Z+AwpyY3Nv27q
zGu/mIdyZGtUpTWzx0MCVL6hKEJKxpz5ODraa0irJal64uUB3SivuPCdWdsqwfBz31V7KiCZklsh
cdGbrNBr+7TYh1QiFZ3BTibpKg9QI2j3xUgVMRq07/hX7yFvM39XW/91KhzMUG+b81iTcdNJsori
mjSMtOYanc3Fk505qaTMp13azrwopstsfkKKv+VZc/wkk7jQ7WqfOmwGqphGJOczppI9PJWo31w5
t/jgINGS1jd32fV2vqV78hZzD8Zd/bt+/kPJMaStivfa3ncWTBe8p6ePNXkVxcQpsk5Y/zTXgNLq
jo8Cyit8xNrzgtyM2zsTUpe0XmrW0Q0sOH/KKW+ZiyjwGlp5OZilsVVgtDE5AVzthm6xKucLCgaV
AGVXk12nuNrE3gdvbvN/Pzy1lgG4fViLby1V98RTHt3ROjUhkaYXXcKQKGwZFK/aWRTj/KaKPSyR
PHBIXdCCXqwJufvo4bd5cHzo6JbdfwDB9+tX4/GN5oHhXBY3VLIsLi0wkQ4YwYoDKEygogWRH9pL
JZxCf3oi6hqv157XSfsQRSA5kOKVU4XD0hY8FxB+zXU3lzMR1xaY6eTbOuL+cPh8K6RYQGolwVXy
R7m5VNioGrklOyodsaSXOCThkfTXKlWz5riozmpgwJJGhSfiXXNbhQPfkqV0ypMW/dtRqrKPCXqe
Hp2GGJDAVhKE0yvWUBGtCTsYINKRA+Y/aW9rOmtLNURfpQpXypN8bBgmubr9UCA+PldjHhJ7X1B3
wfpbzLwrByLBPuZnD7S5pIdt1jehAuW5psxEJZhkmEXjf0YTyou2C+veE668m0wvvByM4bv+MmqM
/K4HO4NDngS7VfGvqbi0l14dBbyWot1C+Rskt+G/QT0Tjn9NBZF/n0s0rbbflAG7zZ+UGooqZtrB
S7Tcu8eBC37lQbuBd2gIsKAbzi5LFg00AkakHBl7mv1KBScBVZoSaoADrGXxBOyR9E9m7Wf7Miot
bLqPT5lU4zG4K0rCM+UT/7JDzY39StnJ+UcETFB1Igs0X3LcSPlvT0bDI0H0DRu4/MQKHH472qHE
o8mkBogrCwQcMF82mb7vE+QJ8aYiN2levBgqavbiDXhP8G6/whBJfqrChnqQQbMecc4z26ulPgxe
TDkz6A4xLblBM4w7epu3Vzu8qS3E2arVkm/Ov83gJNwA17oGOPv3ZwZ2JvthLrnURzyOYwRgSuNP
vLaerazglFoPw4AxUiEUcHWkpHCer0O0Sq+zg3YhTB0sPg5RU4o7qIimbTitxvAXYMj6VCEl0+SV
pWMZfpWQwkm0Rmz4+iqWldKGu+kyF1jLVRvt85Va/fx8cZYQrEkNsyxk7OdElcGwc8qJBmnbGTlK
fWZ53wb/lklUcrh4nEqqXBJV6va4ax+JiRWbRKAp1mZHI//BFU637ooy4IHieg1wydBdxWhgWErb
lGTj6HKKPrMUyKLG2TWxtrEArxSXSCK1tkqfD70Um1uVt6JQlIOEYlUVHsiGoRqpLTX5Y2D+su3S
wut9qjpJM7UL1Be6M77c1GRZzLzzYBfcbpcHyX0zETuNTrMRrf6vqxSHCdZT/vIHQ5UddvxSKhNI
TR+j4TyI6TROAPokXrJpyFL1DcDvoaaMs61enszfUX4Fegu+bIyfEuMOSGWoNT0KPGOo1I64I2ID
XxXkw3ZHvxJE2TrJ0JWQqD3Gra5WOMaKC4BYxrozMV8uWbFjVcpUdEjT7Y5fFu4IgntFkB/DI3+w
TVMlBxBUdUemfmL0uZ5QvvfMnaLfNCZtsGMlfQyWLRb0Xz6PmppR5ek7Hvf9yUcXmQaa0NwcBhOr
P6Z201ZKSyY2NLUW2GXDWk342HjniJQAs2alyVsly2otS1AkrjAakJlrhR8jvToJ5jTA9Alo69Oq
yEKM4P3vTk2OB3bxw2hsOqYtFeA3IFGs8qx83N+Cg7ICwT0i5oz4y4YYUHAoU5VISkXzL1u6B1TD
eGFLVTVOwskdhzjm+3WdDExRaS3u4loYcUdSPJWJL4xl29oIL8CNO2joouKd4Ns3i7nz4FqUIIqe
grW9u29sb99UGrsO8z+29tJJkKlE7pcuCwlz8JObv0x+18NgO5YqpNhFQ1i05E9XIQlVI630Cs3k
zwf8lw3q/hU+53+kctZwDZqDLBCQIttZlD9oNvuy4BA3WAXVb5HLwT432b1Nf0LGeQi0bUWb2G6W
IJVlOWMXNrYuzdTJZw9JoZyEcaUwcD3jOXW5cHo49QfP7FenZ8xQhpE8LmrA+uGgVLcIuRqcIWSk
Uzf36T7R08tCfZT7zrR1r0/KqjM96H4CHNQWOdzhDuV0po9UhzMmfML7sYgHVM47mP85ipnpyMj8
e37tE9sGno1h3arkIecc1Xz7xvyEvja7dfn2ysb9BdZVU4KK9NZi9JneLluVavBYcKIYTShq6t9M
bOrIQtE4h5Q9xaL/t7TAsh8tRxHQkBVnoBBI0HD4AlA/H9Ae98G3713Go2paIS+/SMxvy14Uvr9b
9JDaJyBnGr1WX6Qc7ifNtbLmGtS8zsqm772LIOgxXwaXuE3ERZuFhOCvwhIKiq2EFQ4RCEq/kj/Z
fqm/64e9AhaifR9TPNQFVu5P57x5c+oJLlUa5GqL9ln5t2TR6N5fyETMgceJCNDU8bhQRG39roml
LuxwFRSHzdLjB3+tnQbl4nsWDG81JoS8jD/DFiWA7nP7MhX6Rs3aOupAwyVSSQdVwq3h2mM72CZm
L06hG7+Yz09V1J5W5W7Vh7rBaSpL4PakQcuOJ5XDkKm5r4vev62zADW8xaEFobQZZ6cneY32nEQG
pReS/ruxn8aPCQhVhE5NMPwx58kFcWATePWUyyncUYDSk2NMyjKyQOt+nUnLfEWNzCcJpFDsUGkI
g1dP1tSdr2KJzB8tr5lJu3xZon/kVIMrtSzzBWk5Y7ejCd3usA4OAoJQvnbx3RpOCKRq3tTkWD8z
zc8AlrX4hqzT5MY1a3YZ/AuTygeWrPeD/OZbAEpoNNeDgI+XT9OiGuaRwBuWlYyJnnnaTksuN84a
tz02vsFMdlPg6xqqczCmrYYAOjVpVc35ZdbAdR1VwGrU5UZQnadEn0nzaIgQZ4KBU+KbcjCtNOpC
XbiaaqITGUEaJ/HlcmmwMy+pWbR5R3ucLHQ+Tv7Z/ROAMwzlW0MYgzWlmtnZxoVJDiAKYk4xBe6/
jkBHICezLknLrn/jVTR20YuQCiFT8Yj4LOjEYDZ4rYKgxmjiM6MQIh5I7TKhG+Q8I52kXfYQbkSp
Kt229v6f2l7jx5rgIhoAoWsynmtBytMlQn1xNkV1M6u0T2kUUuQ1sRPLjqiGI2vQk0MqZeD9pzyZ
1D3qEk/gxHuzsOyypRo2f/CbMiFP5U3YAcuNeI/Eov84HHKkw469B/ScTxUqzOeoQT5fjqmF05Ve
oB7+Z9NlXm5+trpSQ+JHDAIkU4h3N4wZd4G4ZWk3PhpiDE+SQfp1dlijZHJguih67CYYE3q6plNp
ZY/CGpfee6/tQxzpDIZZ8MSdu9cyZP48ZAMRgo/LjEW/g5P/VEa6UY0Vb82wY8W4fPTeSq9ifBcd
C1ZgSsBtro3hwPfgmGB6XYapO/q3zkQK4aag1gyxJTVyCc8E/CknPrwmlcduk9HzRTXH3e/40z/l
y3WDGEgCkSBFyp7P13Fm/vESSISN7jqW1jG6oyEkzJTYRf2lqEtvxg1LF/3uAyAMzo03QyrtXkc/
tH7vWsW1T5GjnGXbS37/iWCwS5P6zvhVktyxMYqt5lO9RCptQ9EvQR42EMzSEiatecFk/0cfM2kK
31jR7pf70oUV81nDIq/WQifUoIglI3Zx+3etIgzt1wjO5aHGNJo9+Z5LMHencowjhhVt30giQXHW
LzElBFzZEMRYIZNAHXowltBaoNAx4XxiYt0q+LQSfdLEJiOzhBYJMOKxDlgjuelkstaU1UP6NnVM
zN1QnjlQQKmPH4mabbN2uNJ8RbZiiBimQzduv377ooh+VkfFcgtWoivbtrBOYSsISO2S/pGcJy+1
KU8cZMle/grR5gmlnYw0NtE4LyA/uxt/z+YKBwiX0MMIGo8hYtb+sAz8IqRALiDp2VnwniAXP3M2
FtRh2yhY4Mzr+PEtXnNhY7bD1pB0OxNUjKvErj1PMFvtdYbVH9jBwmNac4kUOg2So+vXJ27Sht0k
7sHPabNlMHadAXyF+BoR5y65EB0HtOfhkx+Rq3pBSXLTfjZrx/QmQyrZSd7l8i5vLUFJlj82vBHc
6G89yixCFYTt9pwrcZcbCw3a29+AkBMVbA9FbEwHDEBBCqtxcS3vGes56EcDirCWF54RgClWhXWh
mKHqZ6pFukna3VwCW2uF0gsN/zV/SjaeGZJCGN0fcjvwLbKduOLOZmW7qAOxazI9IHVxksaWeS9E
vSOaTGu59dx65zAX1IIsPajHvS2rF4gcEl0BtGI0tJazm38Ez5k+d7DFHoqXOwYBOoa3rkCCbmO6
JbJUDq5Mk2IVoRJylErPj4q+2gmUQcukT8YARVN9uQdfOaZ1E+Ht+jU1QVtP1cUBC85qxfVhGDRg
DWDEocJn8r81LL6nnJdYPbXkmLdIgVrTYJG5zTb1pzq/utofLlR1/QNp+frXGuJnJJCCM/czM6jE
IqQhA3qZysBPlMDbqe7RbW6/oyu3cXWJpA/6fu0Rkye41rU5Dr1vJ3ZcNkoIsKjjeqfOeGHkmJsm
Mpi0wfuR9fOGKlK4K1xEFjwFwtzOrc0v/cn0bmzPoLuF9DpD8K4QAqz/d9DzeRZi2WE6OVO38Nxj
VFvy23e6zUK81rScCces3AB2BJbD+lo3nm/Hi18HGsb+3Ul0XrWXXdACyp4f++3s3mP0l+wjJdWP
nyc4wgilFs2495PGSdjFuv/sW2RuIo3TcyEwFcWncrZ4gqMWsk0RI0rxDoVhpr37tdJhXWeZhWmj
Kk4Exo5wMg8Ma8BIz+NVrLx5niJePe95u5bhh6sHgDcmnhCij06Jgk5VhodtO4qqwyzQEGeA0nHZ
Wb6Ye05Wxx8nsH9eDhQfl7St55SstTftY9W7Bn4KDmMSzniF+/pIwDUP2Zucwf/jF705CBwuSCE4
lTbBM58GPkYaz7/CNFHJw4PHnzqyeCzGMdmY6wPC8UHJ6cu4fw3yRSTbpBdWc50UoOfN6E0/TlMp
/l9G5PL0HAdlHki9EHnNFrtMIgUi3pMEU9bvMoItS1XkuP1J8KruWuZny8eehi2FYv5npHz357S/
xtmzLceC4lGUmF/59gpJWMLwzMwXmwJOuj9XHiwsJDKYtN7DbXz6kmN9zqdqzZWIOyDFgKNoqRIW
UmyMnUF6GrJ0sElB2Zg3e8XZL/etNM6W0dWSOA5WSs2veQwoCc+e/uYKNBxrkSyk3dT6xLvJnbpg
gisdvrzaCXR5XeW1f72jVcbb87jB52qlkYCSqFbjgCppNgJ7fdGmYuBLIH5bW6z5AC1w5ocxvUXe
1mlACpD9yx7h9VzepSALC6belU8KD5mfTNyEPgSApMruY4NlzhBXc0S5nhSouF1XYOlwtjZf+cRO
l7ROuEFxPGEM+rLk4FW/bFhc53k8dFpAwneeGWlao8qGyAMmDj0l7IsomOn0y4tBqoDmG617R54j
nukSVYfoV/FdchDH4pXW+1n9JXJkTx9gU5pey7fIW14EVlng7/Or/+162NWTpXTAJs5ulLP0wQT0
515BeZfFd+F0wPy/LQJuaALKbqX94I8l16DuX+MzXpKJcRWKE3PAn6nxIaZXVuimqteA+DBAlXYI
no8KgwHJ0LhnSxlXsuqvS4K61Rj7xakqs7mPI1KDTowg5AfY4XTcBgo4+sCe8GDl38526MKB0nhX
ACuKiJHmH5fMk9Tt/ifYiMn2aPk8X/o3gF3bx8XhVZ7Vp3v2K+R6wzYWvs4o0q8G5gkEfH0djeWh
la1aFrHQtIWygVrT2EUoafoMyxxaalHlukr28kALER47dVex5BGAPNZl4OI2eQd/buPiLvoTGlSt
SGqnWhob/qRbJKOGTfxUg+9I7GUsGUKGxUxNlEnIQG6dh1sn/2tEPocAvfMM5QAgEiasDYVCwGQ/
1nW11wJZJZyImn0k/hFLAld/XNWyxDSDlegALAg0stcJHAWcXUGboELIwa6Tr6hQZX6IrpSfGuR/
zPOO6OXduEZY5wmwaeKjeczLL+C73btOLOF0zV2fXb7WSfBh86i0A3wB5DegIEY4F0hsWuyOSapm
ltOGjXiNWipWwghhmgyzSD75YZ0n9k4AJhDobCqP6tBxq9HkELf8O+q+prSiOxUz9e7qHFLMRG0e
HOW0AlyB2zrYlDpzKlvasMPaZiYZHe+2o3VZG7/Y7kWGwdlL+seeochP6YAziEen0c7IOSfiwHD6
MwMG/7BrT+zUYxO1IlvaRcXpZ8D0PJKv8Llc6GX/pYi4m+vdAXxptG1UmAjm/zJZonTTCvaQ+AJL
3METNzkPyomXXWXMwknnZQy6SHPLbkBb8kZn52m8/tPeG16zQ6c8rh3E+7pDzqDPSsqJ8C9+a4Dj
8K7BbODWSRw2YZEE2n4vg6py7EUMxY0SBt1ExC23zsXJhw5NkMTicyMjdj9YdjF2QAWnppIt8ZF8
+JalQP6o9b4/KxBx2+EZ+H6g4DrPVzPny1x2lMdGOwIguRV/WNS4kGgxBPPWXlvOGS2RDYV43rIt
pkdmZRrB+a/Oq9d/WUqzdC9FNr8KeDh5SE2d3dZ80aa2M2jdVJwZ5wuWiwFI1rbGKizPxnnS/eQn
+BPEZB1xV+zOUJwfrY7h6O3DCjQxUN0KTyhrMAPH7I6acBAZHT4S4fo5Kd1QFxijW3VtRpoq/awu
s/3Zxp9ZtTsc/LrNPyhDB9KLhVhmJ1MHHrDTuncuHhItpGgB9LmBBbhj9N2Yn4q4BwnmSxTazD3R
ERmUK7G1mjNrX+vm88dApfP0QjpfYXVmY4aZ9LFYYrSLWHsYUDPE2vsoIduhf5vlFGXy0m2Tjo88
Qr9W1RKAxGLtSBVVtJeYZ5xySrthGhc/okRJKZpPMX9sL26it4F2LLu+WdC4jB/dHOqwVTZ7iQuC
NCoMkGE+KbSozUKS2xdF4ARzXuFTtI6BLOqJkNZuOI5S5OYBvlU+gAVk7KtELWx1tS20nVieYond
35kGrq0hyrBsD9Oue/W2RxMj/uJp1+KPFu8ahtPZoS8y71+06Su3Clp8HlSSJPMnSvHwxBfjKugz
mFbaWvo++khbY9wuZnoFLdL4X7WA9jCDU5muNNSopX2xxW9AtL8Cijsi2o9sv7+LEnP4itp0xJtG
UiCi76EEJRatmUVlp3eYC28e1LRmED0AGBzz7hnE+B0xSLEd991PUn183fO3vL8TUULUMbejzf23
EAk7mjNcK2gvd04nltftYgayFA4jkluf759wOw8xGnDOA8M8V1x9t3tXXa0wsM3adNp0dLU9wJVJ
xahUxN7NZvdNj21w7Zfor6N6PT9rvADNgffXZuyRaHyz9Kvsirgne+2X6iwHXoL37S7v63lJ+EJy
B2+rdrnb9stHtYimMMK8HHBdRQ2ahuXp56A9UjqhZID2+W/LyB4lznROnocvI1q/D24oKmDfls71
9R5GalEveBNVx2FglQUKRaROBiXOVUpditdcoFGAWx/irNZVjyGNbgdfAG8uz1qUH8nJhV/K+QA8
riVo1UmeA8vUTkYH4/cMr0oxpZyBVFlx53ZgPRUE1Fp4W6wbEiJLCQr5nd0vPkwt54NrWfyu9OHr
VXiV/2eTc5wc6y6Ehp9gA10VGdRhRd5R1AnTh+RDxmtzzbBJejHVlOiB9+1rzBK4gZEezYDgdoof
GIp1J1iyuCQSsaASuo/hN0MozC1CFPXwlHlAv6W8ZIhURnI8lcPkkbut9OKOQ89YCUH6ffLkg/yq
CXSdoKyrAlznpYSjazL9EYEEipSlCLUlZdmnkeewYbVJmCUfTsKT0n5FZTd7vC5WWutj/i7cq6EW
oC4ziqP3hzmnIH+h5uXErLAEipBeDnoBkkD/dwBFTrPOP96af8s456O8slMEyrByQ7al9bLQ5P/i
sm49UjHVwVDkLLAUQUEGAcQX5h1LuzGX3QPeePAHA64+lISi4U6J52pfv9vsHWutuyXVbW4rTT3w
7HWGqoqkA19SC6acMKQbBqwuW7T7zH6L1TahdWipojEW8cahCsSfoSchFcc8xhEu7FW//CSOACbO
tKdy7tNwGYax08U4HEREEiFSQYSBABHODQ8Q2BaW2jsSZgSHbnr4O5e11SZdzivGGxMSBEbVYCX/
xwBtrVlZztCjVZwY/CHfSjOEKIVbzQq1iPq76wjx1KKMcY80gP8Adth+bPoJ6MPliCE1ETNBFzVu
/YUAabCRVcKYfklY3vtqo8ovHHthzEwErfSX3uJMMQbavw2tNcxH374skSM5DtQ8yha8aIrd8Thh
x1HKO/Z5RDJxwj6N7zY9rAlSl5QZUxoQFYYudlwaVseCCuu3/pDzNJYxYblCqs+o9E7Zns77OrM2
DWBCYG7/xT+467PRTESTis69kQKn2KF28M7bf1xDIHC37vxwIBL4zzwhY76wBDazmcAqZWwc3OFe
JmAeJBAWDEYQoj0Ce01oCQCnHD1WBVMVkrC6wzPDDMh0ZmSsIQmpKSH1iGCV4SLk3ThMZlHO+DHB
aMRy0SEUGHR4RFcC/hpG7H9pdK9T+XeZf99JSrTfR7TS3rJzA1D3yrspVQ/ooaRhRQ92UkDhpqPT
oHJYsELktv8JSqysuKrXjCD4l749Fst1gAItMD9GfbZ8pre9eKdUOPrvpTeRqQ2rf9SE4Jn8xRHv
p6rLYWK6X3WzU9vcWnn1nJrlAGoOc13HLnUyH5KhWKn0oDBniquEqC+S7RUWsrLlRqqWdc9JQIVG
N4XNWKlbe4JgtzwK2tjGQydCBx54jzGIi7ELlr/8tZFTF0XcLvl/O1hkW3q1/svfdzoFmi+OPpjl
RBy2vPHZ1bQYZxxvETXPZhjw4Js4XgYCcLf0ZSVQoYGdBMSPDRHdVVpvReIWzV2u+85mj92B6ffV
srNZt6CZ3TXn+WnTFDvQaIc64hFmQD1XRaRb337olcSiSqxfiwdzz7yzUhzXEmYCcW5MWwS89pR6
dpRKOwCUIh/ewJ42xUDudCu33c89InXtePZo9q6+/Hy2DJ893lTlSLWUCXwilTT+JbJjDE6c4BGp
grSuVj5qTkN+QK16FzlKZ6+Zld+V4QXdo4eqUZXAAcrD6KlahEMcqY6w30Fc14Dwcv8Nvz1U+I6j
YLnWKokDdYef64upn+yp+omC3MDod++rIwX3SEoAgItXWKDIMG/9DPlkTTmUyQszXvSBoiqSdrlZ
r6FFf37FjEVWso4JYBKoeWy4+2RLKB0hFgwVTOP2OPzy5Ji/u42AO4gfqmNy3KBJjV5oWyE+lGyg
N3rbdqwB8EMFQlNu7mP8riP+H2VDUWubD6vY8rXCmCC9lvRtyL7K1hc+2gJjstvVFqWLxZfbpnU5
rbSL000Z8oEfiy6NpbZj7Lc27oiD0U4Yz6VgKsrYCF+7oErAflJiXMyiky2TRlhMp3fT3UTTaNoX
4KURgmhyub/IUxDPz8LrfOT0NK96XzcSgf/SrEjZ/xvH75Uw65nLQ1diTEA2mV87bOkbl/uWBtTl
MoWVAQClvUX4yDepedB+j/4kIoUJqkNEZzkJB3j96akho8N3EgGtxw1HhjH5+RVokUMQPqNgPD3c
U90ELRNTD552eoTJ1KC9EJFBL1S+q9ALG4I+J5V9rL5v7+TkpvesOqvH5aeE30en3QtwsH0Gffol
yuVJ7fNxJ2KL//vfFV/D3P0d/10n4X6/G1DWJ4eCHD64+f6Eb47ZG3qa9ObMlcs2AwSm55kHkz1h
mYqR2KxS4KnRvDjnreOilm4eaU4BacQP0JUo9+pYuWAOGnobQsikPTx01g63w8FabUIQvRC2PpAf
hskzXk8em8BFTXxaveFGpMmIxQsqUXo0+x/WuU1y0nEwuk43POXmaszl/5LxL6p8+3vEkwDR2+M5
PUOPmrQI/Ej1RtuUI8KrX6C7/sE2/6UKkvHARZ4pDtvrZpmAB9t8c49Rudqg06Ga7RV6e6aSwlhq
o1jsNhyuA7CWkXjT4BgPn0LVnmpAL/VPy1HtgUmLjY9C9GiJHdq0xbFIZ78Q13rSmzWIUWLHbVGm
7+gAy4cJz9gJaAtUvi55FC+dpz/Zo9WfBZCfX6FOiLv6gRnbfksSHYDA3WfBdCy63I8DatgCtaWx
cyR5sBoezueibECEoUZMT6W1y9Fgk8/DvUX1tM/0EG/xhWtOG8iszCP23cGx+k2cFDmDWwZtj7b8
KAEj23/PrA2a/7Rsw6dCaDTuDyWW3r5jPfpgfXCPghIz51MP2l/9Gmg4cpwSzEzDtwOGpY4mFhjU
1Y8SCrA3Wdt2givc9yOzTA1HmooXR1dUtkwybo9Z3nubFjlWctX5QKWwAbq9L5KejutD2/IZ2geQ
l/1aX1zqIJ+mVK0frrbfOoyoJLFYwllS4hTZKKl+LVqnLeHVM8qVXOKsvxNst+cyonw7GbQSEylW
gJz5Z8kGgO0JwySkXaC4wqyf3J/HAdpDHV4/bz4r7mrkQpxJL+yIdOEknOJmKbm0zzjoUTuHiUhy
RIGy9NJU+95ELpJiP93PgcdWYG5G8pfFZWiX2+VaS0KlMwVTLsWLNOi7eYkj3uqnTsOx+OZb6jOO
OWcTgN9U/39hHoxMh25UOKl66IL72aS0/xl1xXwm5sPjFvKLTpHYtWY8fmGfIeuu54FXNBQO6Yt/
rn6nH+jsHLARVgSEiB3Fx2HYbzfaBDKH35RewKq4exyv9kus/XavGQxoLvSte79yrrZ0rV9Xvgef
1cPct+vAAEv7gagpGE2ZikZK5yjYI4pNyyk8x2npTtzQS6LyAkB7Ws0CW2U/j+2kAc0RngwPO0s5
0PP6VpEHzBlVOhr6Rya0j7tdJrVJCWTlRsPZV/0NyAm4pEloj2y97MxSjeTNEIWUg2LvHLJHP3hm
RbwQGZaExbdg4uK2aLmPRM7jRQr0WQO9LcPu+y3F2ck3APY2NmfO48G1aDosbo2qhflyW0RV6ORE
mQNatw5QHzoc417nxB0OOhCBSqtuUS2A515B2xMGAWgOqelhKJQ1V7yse53jBgGo7LAETPdyRCxh
DP55SihLCZUvsc2vB6b6Z4BnvOMLGxJsf2gyd7hgrJeqff9cQ6c+QLy+hmjpxgA6tGN36z7rNTRQ
qrOoKlJ3OAbppWhKYQQfKxuNj0xEgNwnKXUgG0bDJbM3vx6rnZnH6ByCLvyCOWyWGtJcP+CCB+Xm
mgPLIEBCZAShIikViqkkwGhBrF/1tQVY/MS0pLE8sZT9Q6JdbxqKL/pSzKWh2UL6xb3jpYbJ4vzu
IDjno8KerSwZRTp2qxloo/O+dOv1dRRODA6aXE2OWqFAk3BkKOvhDjnjnOBjPwAMmZUL4+n6BkXD
rVeKZvFJvg6ohG956zHITP6G/q0CLdccUu/8HOpCugSDKpGq8+D2Px+uv/U+cGILIa8PBc70gYn9
Wi2+1AgCla/xMhKUniLZEAdEb8LtkljBFgLXr34lv3lE0NGb54TiDlMMA/6Vn26W2+gJBbGMDePV
V0go6fSV0JW2MvZBE4iz7QdS+Mh+mJx9B7cI9l4om/+TJwDdzX2z1FKfV4p+e2C7a6qbImIb0nO7
6c9AprfOiT3IgD2Fg2htIjG7Wtgkubi1raxq/6EFfR3W1iHwqpuhiUmc96QrXqsdEE3BrWobmP5T
9+HeH1pqzRAbw7/lu/pAc8c+gqifGK2NXAJBwhqzZsDa5912nC1+c30/5OKSCLal7tCe8/5ePFgq
FPZ3rBGpvw9NkbZW73ash+2eDSI8SFJxD1M/bLV3hXhgW4rfpn2kyP+68NF9kQ8N+5nfBFd8/2oj
HJqsiLR0RyZP0jQh6jpVGlK9PuXR8ExrBEdWVEwARchbEBQOj7fiyFLN/V4diMeeW/6o4048AssX
1409yDM4dX37yBYporkW1eyh8kXCAnjuUzqrqx2AKFVAxa/FGZq9fRNd53Eu1WnB/Rx+A97WJvan
HPwSVaMql1y9f96V92Kz3x2JwkQLFJ7X9kuJwoB0nMaH9PGIlAQE4rOQf9PXuDV/4S/LCnizFEsX
fqvo0J3BwSKSGxbMmYGLLlw7hL1rx0Ql+MrWbXK2cwPrHiZwtQUZXrq9QtdNWo1gJbDN7TrqdcDW
uQjvS0GsqfrD9DJONIuKIO7xrrJv+aC1jQbGANt+Zktlv3jKyg/t4zM2zF3j68W9w2iYp9S/BIRM
qPDtwaL/VnGOfDGeDQCZrYfrlCNLqifiGguxmL5yfhegw3t6Xf8nv5QIhaqZpQoUMNv3/RGBixyq
O0Kt2f6ycSL4zFlQU2U+wX5U6bj8EckPZ5kTbkkhx6Et5OOWVcWlgPRj1wwCyQpJD4bH6crRijP9
NBVBELySZSlJxR1XZP2eMOcqtZkVtd2P+fHmLzaCyUaRRLjqS6ViXMrAcmLruw+TgexPj7sKU8EE
HJng8NwZu1h1wR3MvHWU+NOX0gVpJrDTSMMLr+ioNJwVxmVGQPq9CQ+hhxOHL6pXzXgLX0e0+3R4
gxclG3/+n9Wcs+zlmciefAD0iqx7c/BHkaA7iTVGaecr57DSkkXUiBAuJq+9mL/4zr6y781mzqzY
K3EP9iTfe3YhL5N1Gv+AMSjmh2h5EjUH8TstIP68NCmuMcB3Wjmx5WnVvDlMMubwfeKY5yc7/R8N
jpyAQd1CtsgH0S+2KUvpTtSisGPNracNAZu+dZGXdIK0sFEvP9VsCgfCcBvKpB19lsuxQZGrCqZz
uJtp+tCRid6fwZfuhZ4s5EXqCaZ5fxZypTlaeXQKYtYurODDkjwP7NZFMvu+3sG6MMeYnLg7uC8t
NmTqhXKJ6/H83ilOTZIBccgqvUrLE++IMgjd23WN5Rhk3g9iTXzFLFnKluOtbtDIKnJ6AVFX7Mqw
o7BYiPQJG+vR7ORTC+tAeV1Wn9S/A+K6Pgs4x8Q5mDFOatWKGS9bZvglve3Wh4huxTrMMWsk/G0Z
9nf0Ld3VxihSK3xxDg0lFofCMHdOkuWH3goj6I1aWo7TPhuJOusdoLDh42dE8JbIKKk0zghIVXlO
LxmLWkbqj7KEuS0trpRbRLwEyKfmCoetXq2minxQwzf9CaGhb9ZbKQ9DuSlCwkO7ucZzsEeXhH7s
fNWxEztZt8uYXPPeaVm6OjSO5GyyHpfK+Evk5zomJoRbBldgmv5q7isdKL7Smpo/9ap1VJzO1Nr4
5hiRDnSrWo19htkPirBUMLiVapwKkt63fJHj/Y129j0cTtU7EHTHZStWxppSAmKJBII7i3Pb+ErT
xmen5rdTpjHHH1CNQFe7OiAaLx8mD11IymWjMwcY5L7v8YeGJQLkSyiercNftyBuufDHM+/lJBY3
dBTb66BoL/fkzozfRmPBCmLX6WqBpOV71JXHDmDg7Oeg5uoHNwD5paDAG1Odjql75XlqIUtg/YlY
Hr6Jzk/QvuHdBPd+N48SJg51WCY43jWPlsfnQxcHtDen1KzCxLDmIKQglwUzZ7/Ask33TadM7nsL
c8Oqn/RVh3uc/2Z2Q9g4aU8O/4s36Z9Mvxk0XbAY/HjLgFzgOYLPaPCQ+z5lfGgkrXKv5O8UFdyw
thgYjgTflubOyLm6ydeAHcX7Fjf9cKUMnnqnGHNsq5gA8sR/2LBHlbWP12vjX7QZiG/QbAmF27E5
j08zD84S0cnC8AQzki2R+/Ed6nM/cp2PMC/EKKj3H0aJC8uTqSj81zAV13iNW6hpAnSMcU/K59sf
gTF/pCe/YaqH39BOsmpVqaZJ5gqTq+CYLt4tS5sOCwsL+L5vUZj3HKve0WSnfEJx8kIi5+/dI72u
yF59v96YWC/iMAXmpb2qg49We/ZxlePnFFOLjFneOBnpDzQddtPvPqOZsUOFjh08Tjltv7vy89OL
EHS6++pXVaTViex6/Y4SrERMMfzPAqXd8UKUKytvKjiBlIGFAOoi1c6t2ToFDb4gbC2fTJBzGIj4
SOJmYEFVNbggsCU+X4yyL8ae4f7eJuVwQAlvKnYqOR1xe0TXGKNFhdlgqPoQxvUiHeMkGQ/v1zdb
A/zR4s6qHRBn0tNECSkBT2MRkknUeUkmfV10W7a3Lbw1vVPZpEwC50yEavjhniLiLha5jveQLI8j
BfpoWnoT+/5cghs9K4dZR4iPH21Z8Af2C9btwffhTWyQr9yuOhUpnngaScEoMY9Au1xR7ZanKQ8O
zTzfdZtPTlzcsHcNCBYR4ygvXxDwV0djLulPFBkBPAJEKx/4F+o1Wcd9QAqvwbrilXfxJpznUP88
RcaSt+HYC5+VBvFdMVkUS1yCAVpxDzctpYb85aHVdlQ4CVcuhbun5Spl0L8f6a/1myfW3BjQ6YPf
b8AWa1MnApteMdx3BtXvuY2NFocelTJWum0OCJSlvIjO0EafmiPdR9Uscdh2ne1UvoafnrknUuji
F9zMG9qqBNQvvowuvJJWBi/1jR2/Kzlt0RNCncTLrGJb2WexWDpMPiznfGqPQOlp3jDKpizlWb13
IsCo0ha3XPQb+MAVtFC8WLzZyyXKq5Yw5q9sUX3wNgfxiRQ28V9n2JN/XxGVZ9CZXuCi++awKu/S
ZuAnwf6OvXPAqP137w2hQtFOt1dGg0dieZnYx9bytcu68mev3Bn0tp/DtTSexuSnPtRXZLruBWJA
1cJqzAUEpl6tN0uwtlZo2aE8bJ3uiJCotOS+CEBMuBHP3ouRG/Xv1Xz3cmur0GBygS84fvvjFU7j
GUMRB/HE8geqi7KY+k+YD0iUPULMoh+JpzuQorsNwr+N5VEa9ic/DvLVUNt59jm8ou0ZlM02d14R
ADCH7BUse0E3TbJYYi9OV5XMGcahOGFBl0oayBygB1I//MutkBmVHawJAA1L7zJmApVyI13Ew4t0
skCTJcL4ocsZEmMA31kvFoodAU3SpVJZoTMBQGXZ+7QcMmzVpdO4NyzhjJK1+DZrs8oAu3oh6nXv
wsD7iDuHkVD/DCqS7O391OgcOnwFcFGrIQImb2l2SshG/uNOGtsg6cU7AzspAat7gAHJ434fGw9N
kHc7ZcBzM1X/DD2YRzGXWcUyXwPbTxLC8QcU4HBGvzS+YlFM5dDd/PIn1n6gAnHYyGW9iEdhw5Bk
cArbHTivu3cSyiTQrHVPeJ1Mks/jmHB16Kbh7RMDxh+PeMbEt5AR5hXiLGObmgITjoHy+VICq31R
DekaNbpHEvTnFagCOu+m5C47YvaI65i8fk/RRv62BUk242rGMfFWnkvWMcr5BFwgGhuqJDhccAm0
HjmTgNS6DH+OMXNITXsm90n6VuPeWeX3yz/adqsFlaQ9L/eeH0YiiPOAdrSkakmiSpk6/6GkFD6/
z/k0uZx8gUozSg9QJKTzRMsWIX5+o/KupluMFtSZ3eTa7dd1y6DiH74ESOQCMttoyp1amVLBULd5
XRxNO8UFic0KFxIDoA7qMcx69t0ukP7VZGZsYub8e+hDzrAo+wjiXKI1LjMHR0r50a9YIc1ZoJmR
pZIDKykgXEe+C/yINvQQReVy07i7r/WJxDvAj9iDSEZvIAB5IJWk3NhzHEB6rAwrUtq8M/+ULSWV
JtA190CcBTU2I1q8xpgai+NQlB5jaeNjMUB7Z20wuihN2j9UXJxdtB48UE9BrjUAS71NuhVIyD7k
fuZbokVDRohBlXvTj3a2ZEKW80i3+HwBnbjy32cCAevsiVAhNYvz7ub+00Lvwfns2EEoBW+VVXSr
7FpmntuiEJlSPl9bqWubqotSLa+rsJhRrbmnX8L22LXZnqs3+d35xwc8DaIoMhcHSIBFQcU7V71G
uznEq8v+o7TrKmsKQFJ+7RztaBVwB72vIPr/Ek1r2g7jEymejQmwfcnBtfcYJK4DX4/OYboPes40
hTzRR7/s9+08l4PyvbUIEG2Exe2Mk2OSfputXmdy/HhAq+4x+v/D0FtjnVLQsHq+4hhFZc4JB3su
NziBRAtWRZewZ7yaUPwklWW8uDO2Jp6BtF6npJOvEZRr1mDmdNevPvzHG7xWwHDpO1n9FOo05prW
/GTyiezp+5mRAeN3OzvGAEP7anvYb/B5ghWG6YvQXVWlxJ6rDw5CISUwnz0B56oVUlX407BUnLtA
9qMrLEGPstpv0Y6imXyF1I/gkDICe3Ch541B63FcMflDU8I/kb7xc3yuY5OHbNWKfZh0ZGEDgu+r
UavUaPjXvhGVDxKcCFl6ip6J9JHxWWEW/lJEPPt4hEMIBI0SLjMSH0dhbtcF0fr6sSRSFf+ZEu5T
eY7j89ur1b3Akso42nngpp35lny5JqsEgxIfqSZPCuV7CyYE3W5SVQbwKP7vTXXEzVvvUjIeCLJN
689kyXStjYj0foRyJlvTrU8ifT5/PctPEJVKayvqni1zrURviqeCfsF1gDYqFmWDo/a0YOgiSNF4
HfU30nQngo6B6l62E3HLd2+sMHdTvgykLXP+CaloCn+70KckULOERWM/PCIzlBgvElSdlnQLKFdf
UcJe1IJcmMNuz1TJHZKDWWvL1VhlLjjj9NlkTE21Y7Q/lZp+Hm/BHNMNsDqxfFgpTIuAq+WmKSUl
UtRCIf2UPn/d2siLtSKbGWX4mUzMx+r1YhjXa3oxZdg64sMxtFCQp7glu4kc0OkV3QHEwLRNOvTf
DNIaIdvkJmVGBTYLvoWzOWvfkv9zMDelr6VoRYcc9K2O0do8KNRH460WgMfxheWnJzqGLSPVCB/+
lhtfk2HFD43lPL9fca+sC9IRTOIL04LjxKfPT0ZxxsD5ih+mx0MS+mwRmCCaHw7WW9AcCeIcrkh/
sJCAfdGYWl1UbudBa70BopkmHffCh06T+HtE8YQEN9VRgUwa4TD5mq1K5NvCxcjEbLb0FnCbfbvr
swEQeHLFLCJuykg7lxXkJvb3ChZsHpxka8T3M8kjK7uaulcisTBWrMQEa1i/S7ZGFyTttvYNjoc3
SApys7KNKicxVuPqdcdZrJli7lhLuwnQTtggnF49Cub5+/WSIIe/8U3lUjcP4uE2iq79RjLJZvvQ
a67CDP2j0/Iw91bCX9APqiM43+xWXYiP9Q0CRWUIDwZSM/iMHjPfMzYuOQO6cmzTaR9QFRDN7VVM
IDlquLFZ1pcW7ML0AmlUdIw/84t0jJeXFHoYjf1Ta9NG8hYx+AnB97HSzqsuD4ZG/Zcq//ad3A38
ZQ7iRQoTIpzRFrf33Y6QthDjPOO0RX9q4/EpDp/S+sBNZlnVg39Halsw/HSiC6q2zl7hwD6AaJwD
yQWxHTMFB68iSC2ThX2X34lthbu7bnbMYBxh6siWnxnuTpVEmD/Qc3RsxH6hnxhGBEOFQOymHbLD
sJnmyYCaUpnS1aCZXSXd+867D8VGmqJfuvdv6Q2t2AOc2qc+2HmKwsApAejDkuxbUGvRJdB/2QCG
jRPuoCCLR8fGMXmqCnKrYSsSWAtqNc+alpF7y8v2MtDGeeojvrFUNJY9hcpqMePK4PS3EtBTqWUh
LGJ9AjYJy37tjQdT3T3AMzPFY2doJBA7HD+caJZB+jcP++2M2zFauRdmZdpK/QTsPbe1jolRKHSb
YPzh6MtCmSeEO6iL3Hd/mGtv5gdzxw6QWoG4dkTwSoB3Xsf8UOTVxVO+H+litU7H8GDSJuZXevhp
wdo5DIMbxJ2i2n86+feBW23z0pnMh38VOX8ecr8mtEYVDussYJQTaRuQxkKufu3qyWFbaxTEnBkl
yEglffDgRVJWPpz/+VkrD+zEdm9NZHd7iP67/5Ox8xBHjIIcQuEnvhq7wSVGl+TZ1DXJe8SFfC5B
FBwk3xD8Su0WFSZVRP5CX5b5XX9RbE7dlyUAUd6LO87DEezhuY79PoADpC0P1OOTObdmcKNbQTzS
FIxcG/75RrztC87rYR7R3O3P0Z4++76osWqsHCMBAV/lT9uNk5vSoG5X4w8Vcot//xr3sztw2lWp
uAfSvIr5ABqeVPwcmOl1SrEvgpca728A1exLSo+Kz0b6Rcha8B+DPyPhzhHm9GmywYcpsP2tMUm3
HfvtqrF7wfknHXz3uoBt9lZy2yhcM80I1tP/wyjqNI5jDabX/PTJXqs3NfmyxIwyFALjUPfhhL9D
icOJ+cusiL53tlOKgAgq3ZWmEHWnNWfAAm1+RSSQd+P1bquxk0F/fgKi0IN5Qd53pH4T1Rr3dOir
c32atnyAkAkgVDQSF2DU5m1vbIRWkd5Zm7+plqUwCIOISKIAqL3QWXW0ycmd1wQxTBcD5U6WSVZK
RB1v/QtBnFjFCl0XqCor9wbpNeGVHaIiB2GiYXXMssaQoYP8S79wWpkRKunm2pbSAsBULKpyl4+8
nybIPhayr6U8oW0QiALYxLXXuGh1EcPVWE3qUtu77jNyWXX3OEzRkHbt69cfQEGesBMaQX2z1HCe
ZOouBJPlyoOLOM+dB/4K+3WJx59vvbdemHg58ng0iRae7EbasvuGeKZ0kTXq7hBLw57+4qh5JAmz
ne9AtF7LYCOgv8MDLOP1cxgiNu6KwUk/ezu4UIQlq8twaBGuyBgVN/cRI2XY960JL7affrTy9hT9
muxxlqlsbR3FfleZFBXrFwNhnS+3mcfS0n6yeCoojktyczWFIhkB/xETAa0Q3yvG14rlVCD191MD
0gLEWxs3BzpGfh9Shh1CFgbdbOvROMmChC1q1MDZOA+l5X90IORjBtWhO3h4AAfD0maII0sSrvnh
IhxrgEH+sGcOsgwr4s4llYQbwRvytEmvebpPveRVoYk5XNFwStlZZs9MncJt5oMhi7Bd6yi8pLA0
19d9hG/8kYLLlpLJiDeA+1F71ProJ2Cb043o0VEpaMq/BYI2IXKvPZCgKCWJV4jsbuPVtdBTmmuO
ZmifRmhpbj23W/0/GiVkgNK8/JbC3SVZf5cqSvhJETtqGC5l/t368sqoYe2EaxPujhUDNY9kri4/
Mskr3NuxZShV4PYiHbbrNCBsURsm1bp9xfwccXESs3Pz8daASqjs7szSJCoGf2SQFiyKeApbkVC0
mfk0nCUFLnunkXHs/DaXvUi57gROGmkmAtrSO6ZTawl06y73rmiE6O2QNAIDUN5lXnbfU4ORL3CW
JtELsyq8bfxEaDbYskHphrKC87/XAb+O7TUUVdgUsW0YopcNP+y7pCOQHJTe6GIJ7iPLtyz5wDIf
usFAMl3DlTpCbbq2g0zWQyKedKt61fB5AayicjQDjUk8bNkeriskzxFkoU05mOIDbj9ek6tj9b3r
ijS9xjdZMSryNfjaIAi1pyR1YyW6tiw9tNucQeEFAgruXbp99kevO4fUP4Ga/JjYpo0UclKR+bGr
k1xd5YjrH5iZSwhne2r9Xm2k4UF1OAQpLjjCEvbMkpXgJJwIJCQQdPsBoDpKNmoZJEQOL40g1fFn
/hzYzohrR9ZnuQV5iu+pQoOizBmR4TsOzqqNaLhNqGiygAimtyX2gxeyTotHHWVwb7O5nesDyCDr
0Ov829K8FDStFXJPTqQtiVyW9/C3JsaUfM4kzcoHxzW+ah/+yHigEs3F1Oo8h3k/zNc/FoPJdLKE
n6GbVIXoU1Bjhg3mzAV1Bz3o2sfSECPNl5Ktk0jcDrhPpRBCCluJmiWqwa21mkVN8gYYwF+whIQJ
cxjEgLBcTOwd1Ks09x2W+kEk8fBtHjRbc3bGPgfaZUx4fueWRsbztvTU+SK1OKLjK2T1Mwa/aJeK
cwvKUKrcXBD2p+wk/V1Ut68/HiK0ROH2lXc4BRMw/rSa9RtGkDebrxAP1OOBjpHLy4apCZp8+nca
ZaBBB6TuIlx0VCy9L+vaxin0fwgYxa0DYPlPvlxS8bxl6DTMc9iKxUgyoS/lFSnH97gxFCsQpbAp
rPJKYiGEYikapxocm5A6MoKfAq8XdgSjAS3eWr9XVcLRbBB+V1GCUwDutPouqTexU0jV9ly50MEn
yNsN5rmTc3bgsIDYK6xy22n06TWgG+Kte5SH91TIE1trEK9Uuxt1g4Wf6wNoFHedwUi04DeQpXra
96zp5tq9uIu8AA30o2W9hqIkKin6Is3ktXnnFVzGay8QMS+Z5xIUfAMMv5z0oKeSGUVqtwd5tMnn
MuOm3cpHD5yMuJyDDZHmIgLj59+Xhm3QfDkFTjm6va0Sh69dUxO9AcNagkK1ou6tNnDoasCW09iZ
Kkx+A3biisx+0es/Kbm83XvbLOI9cgyviW+n9p92pgMKH5YHCqy4QAvAU65FMLNkom7TlsMCTNO2
KTBVqvZO+GpRwQrg/vKcK+Ubqt2l5YuSW5ZWDu3Bl1GRHYzBs3tpaDWIEX46igUvnAIj8HqTsCvc
yHlCKyQraHqef5KT7pzM4dCEOj+5fFABvxb4/yrr+CjuCU0RikNjQP0koV/C+p3MPyaP/GHX7acS
dmzqyOcsXC8e5zJdXrOWKapubQhAUyGxqcv8/23pJvB8InWnPfl/kBcBQnr0ZJOmN24fucCwzFd1
QZetC8ZKzu6HwjkYc9UmKdAUQA6QKou/kZ9ccwMm5flgH0Eurm7B8zLtSUKz/9GvWRr43jqy9iP/
zfUAPz6DOyrVAp7NMWx9Ki6yyYRM5dfozPqLej3qUipOjZb9YAUu9zX5zbwEN8/ErPlHIGvpDMp+
AYR9WCyGVdqdOVp7SdbQyqoZfX1TP+CWuM+hle66SAHN0EAh+/X7ZYPKwZWUYslfLzHNRKe6fIPl
chJfO2dYd7QL7ssGhD8ie7QStV25BREAEDVRjyQBiTRD2LmmlGNhfuB2c5QSjqkxk9n2QDONxQ+c
jXnv++TaLpUhPaE5fNib1/se1ieZ94dBdCnmBeK8oS6VsDyCLZMIMvQNGzXVXh8prgljAu1kOW9d
6jpwcTmosSBk1R9uMu9xT0ak8dze1H2BQ13bDzrXRiNLWOGp9xh9tbfLBoCkPF+RJwLsblfw8+vW
RBb3c1nU1J2m+oJoSNKc6fhV0TtpLjGqJXosPiaQNfswyNs57HDLg5Ghwmacgvkf88cydtPJofJ4
hh3w3np8u3LYWN1PiMN/Y1JccmMqiz1BfW0vQTAwCvMzNMxVCbOKvgEw1Fs7dQoyx7v7y2fOPl1I
Vt27/h7buZhj3RMyTiRuKPDzUatTvGwxhn8I6I0KsKhoAVdBG+/oEy9h4QQ82MfslCWIzK+YMzLn
t8KXWY0YRD9jWaF+vgRl51cqVzMcDATs2AgwqkNAA9wrBQTpRjR55dsve8uAKqiFdgOGEhO8FVG8
/th0mm9oGvkDASKZUC/ZjVhCFAJICqVmHQII63zlyT3sORo45nmpfhLTnIpWEUE1lzTtvvB6odbB
TV5aDpUpeUbew37fP2P1oRB9mjW55giEykQ0R0z0DnYHgt35bE2cAaqgSmR0MiLatUNNA5GoK3Gt
DNIs24WZA36KeVXmnF0pgrbkYsRsQmu9XNaUl4HlDM4cwqn/5BaHdVf1tj8SH1k4ISExFzUwSuVD
pzotRd++2YfnOwrYdWJpkAGC+8OEtthYTHIz3zNWin2A/Dq+qINJb2v5SB6qgeUiELyazWaQScnW
Jr0xA9yQ7192i82Z0jZh3pCIEFk0iz3UVopuy1X+aX0H8G39/vAab+TOauXh/giPcrOLu+Apxzg4
xqoTZTYh/mpwBYEbxCONDKdhTO7uxIlzCZHp89IGnDokIrG3As7aZTLRYyxI8ni5CjzZIdcQfAWg
QYMYldahy65iFuFmoA/uud77encUSgdqxIpxELEUDEqoSwgxHRVZPgeFDgSP1YFtNwEoQ5hJaZ00
Dxf55PGCaZHYTv5ilP1f232YImUCJZ2WHryQNK3asrEcNlp0K9o3XYmq6TE3OpwnaQ/NQIzX0VTc
eeGYI37+V2Qqwhl4gmOTaAvXindZrLDcWI2NOEyyZ9u6U4JgUR+T4VhLfyjMkbuKnCt+i0FlTlPX
9cKTJGgzjQVI2A9AMBX5yfqNOoMj06XVmwl7duxC3ogiRzq1itDuw4nmCH7v3fZGBOlggbLDqWcI
+gjlNt/4WoFtdAuA7oybpfHGPx1KyBbAtZaplJzGxDSOpqY071NdhMDO+ts347W90llxzlktZ8MU
sjc17GizYuFVHdgBZxlvJBNqAWvRH9UHtZVtr75sPEansFAhW37+uKljjuHUUO1timIp3X8W1xBj
S0fAGuWYcYH99/SLJ0ea41RMmlYkMysKCC6K4ykDBkYC442AoSfPINR8PqZ/rjdgjQ3oX7R9N1d8
sWzw7Fzko3AklxkT0/2aZCiziShcSA0DpiobLPxbJMcG/1LPKMlNLnx3qmNOMS4OkQUhuYHNwJfV
AZOqR3GPjLiS4LmbjD+z8fW7/q5dXQPsRDGpNcUAWwY4QJ4YJXZhRjbShQAjWlNM7YvvY+2GkAUl
FTf/aFEwauE/VvVh2dKpV4NTSLoelzmnECwH4RSiACViqswS7TTM3oHpVz49BTX8nJn2lm727pDR
7vsb6G0h3aP8USZ2VXgtaHp6jjzM1q1E1TnIiTvMIgnKlmQU3JwCUKrWFChVn5ikkeFhYqLhPqL+
gdD3g1jadsHdQ4FLxOPFdNZw3FqyzjaIi78SS+efH0YBy3bNEoasr1bkG9D7bt8WIqbKcZdaSDKj
Amw5lDrqJa5rTNKk9bGOMvK6VjwhC6oNbuaJf4hT3I0DwwVvRoBoFWreN/o6nh2yHcerQ9MJVDLh
Od1QvMQd2HDds9W3tJD11m5BRw06zl6ruXeIo+EegnJvQyECuxDL/EOI5toeaTvryq8uFd5RSi8x
TOz/S641DipbYbl+nBnU1TnJOCJzQ8fi9+8KF2Kwt7RoYSpSBjP+Q/afHvB/v053FZ1H+704TQUu
CaHq70xq6RN+bUoS2hgllnVy0tfrOwEDa6KzBXwxc26KTmoVTnbXYgtdFcQRCom8iBRKp1heSfGC
f8lPixoawC3LTPP/kmeozvbbhSrbW/YRgVnOTA0SwHCVfwq2TuGhdndXgq5izlsNnWRe1VZEszy8
GBN0vqks2r3evVzH+EUMguPLMHc5eIbSd4RVXePMSsNLylIhX5jr6iG+Gt0SfJdrTJSBF2W4KgXT
o2/dgCqd4tVcfsksVLhBR8LBE6wyhmuOdc0eBCGR9mzNDJEJ8mCQnZTAMkU3z5V/HNEVgHU15w0s
BN5fXiwKk4Qi2dw1yZt2oTqw4vBkQJ+uhT+JE772BmubIgoYhVB9dEIS5aCavF0mzMBI22POZaT/
gcIgZXbIkbdUKnF64XgW2zto7aOxIqE1DQrutF2fJZNXUx9Ou0tPBiGBluCa6Un09MuIW80KX5gV
PFK5wOUEFqlzOflwGpEIA4j+opBdfSX3qJYWwz6964roEfj06qoxh9WatlPrIlRBZjb6bBP5OyYT
/9gFwF5uc/so6LN29qvGK4pvIPXjK1ijUYjNrJ+4ijjx1tCZnnWHzHa8EYWzHyiqQogyxKVsCZAz
tPut32G7toZnoTtY5CMn9ax9gl7uEbjL3Y8IlpPbqiXJUq2lrMMrSd7Y4Ka1JhxWnS+o8a42KChC
Nztx0p6A0bcotV4Y8l7IX/rDsW2AO+XT4pQ28s1KU0JSdBABPO7riIug2SSj8JbdxajWI40CEG9k
pWH5/QgmdTIOMqbGzww7VqU4TN2hjWH57kS9gFahdHBQ5aLxC/Ut5ttk47WdfbTxXH85hOQhc7FG
hj9uv4TiMBXDMaVIwgNKMdZKuHbE8vDoOrHGBfT+Y3ehveoAYNMXrbwgwAD+uWXpg+owSV0LRaA9
9YygfCjk8rK22efn1pxikNPi1ygbxrfblb6wOdc324H1aKE4BLN8x5OsBY3ml3/4IWqrkHNCLost
AM9JEhu/l3yfjIEs4xp8Iz2UoxwRLbkP01tqCbaAFCkwMnlAhD1MLujv1BhtJD2+vXgV6kraZNqK
iIdp8rZWSJkI491KXKTzx00D5hsvf6cPV8NT4KzQDgQjPQb6NNcPf9URPeBWD1AlbJzZrFk7kwCG
P0kuHSCD4zpXUb2GrqiPmkVOXkR2glMbiLYmDPJtmu+5YMF/jBKNynjnth51XEqbTBXgVWes3agN
Mfh13S+Fx9SvQ24n2zn4CvkInsnEyp2qrGsExsL3vewOBcUVncUrgoS3UuslvubIzaeieobskqx6
i6XdhHZTu7o4TMSeNGw0TUTpLjd8L79/fxyYL59j6QqxqKBIty966EdpFhrYf9z1CvZwIZD3kfNH
aDJcalWAAc6qdaLRTFwKirJKstaNVdLV0h2ORv2qMrc1XXVSGIgwXDi7w1uWOzS5WhHYaKNHm8O7
1bXlCY8/HNidRs/h75FfMHlD86BeJPV6UtucijBMD84dYW3GMTFkRPdfiGH0AFQJkTvkoGwPFpW+
xN3p4gR8jC0/jpLcG6FKRf3qNueRu8yrbW1gNUgQ6XTsK3sbmqeDTpAI2PhslIZBkwE+InS5KUnV
nLoaxBKPEn9ONd2KYmyG6Ak/LgKZ6h5IaYDhV4DbZyw2RzfpLVPLQf2wsW0q7msfMSQDFZzbl5P2
PYSKgGlIauv+sFF1Dy32m/aMAxKu+k8Zf8xp+l7oPXrKn9z8ya68of9qomuTthCUetpGbEbfwQ9r
/f64rWRf9IxLyUgy6uKnlVHvCgTgTP/BcDc+c6k2TnWw957x/hES60rsnNKOw3eIMdSOPz7WNy91
XtPDBS22neskjLB78TkMXNFbCriUyrIh7hctbSrZHJ5hmTU1xpS0MiG/BWutGMtpXZAt69IwRhwn
qS+qMyTHpy0FARFv6wNY/Xb0RdgOYeGadjuuJgiMLqUSS/aG/wO+GPl7yAh2JyyaiqNmRAIGjGRj
5GMLiTikkBOnJCVDhDjhn3hK2Iz/Ei6Tz+R5dNOI05D1TJ8/x/r/WLZhxgMWGoeAVKFO6/wFdQxO
LHlyICCPfDTFH0VZ1tUWQMzvVdiRrETF4KTLwrfO5qiAExU0QMTw29PFO2GmezTZjTT9Tyum+sB9
+unPqBHnmnCbGTsYRVTcsGtSdnl3/yrBrEyOjeLic1G/PN3vxxsHhEWrme+GtpDop9F9/NWOmmH1
dT6VfY4UClfbWC+RqC2jjCnalWFMGQTCaO2F0MAJXNAVxxggS3YkRJ46f9SPoyEkCdxkjzUZdU0a
CGxI+cNU2eOeuh8RqZUShcQLw/azlD0BQK3MWQ8rNA+kHzzLzsa4fe9uGM0vzadDfS9ltBRFlrEI
tNhCHU//fKJBzrZkFmSq3nuIPBQWtLTH2pWhJzYuZRe9ROBIaSkjidVgzKEw0uBqrVHTosJ5e+bo
U3US1+nBwZAipo9DcuUiEyb6CYk8G/9/cDMOSXPQfUhkOrVxpgdQUrxo82PlXW+XHZkp3NF58SAP
OMcIRsBvYnva27Stv60SW8jzu8slLBFXsW8SnWBtrCLQGTYdmCMd+8lOJEDkbsEcpV+4uEd/20Cu
BclY84fxEt8/cjbd//T2DDdFDhQTeZxIeNARU+hJQ3epdWu/EpLY9m8ZZenGvsjPbzHrQIv7+8pW
5+Ciz7sOeIVPovZQSyyaUQWo1vRLVwdIjMsHh0yCb/rbLrrnQ2RyZpUj1dBBy7iD1YbSM82uw39r
P/sOXyiN2XbGvV7PwvEqd9LTfKYGbihaXvLYm1rv/SaOvuJ6au0Wrr7QfjFlTzpcExAI9JAz/zy9
ZGR2p0NWNo72X1uUuaTzT5EV4JowSGpdJKmv/xQt3CIPDbsdNLtO/TooFJX3sf3lbq5eOUn6BEn9
SszxvtZ50rJEY0SMq/Z1Pm52ST35LzcvBImjgBNFFEqlds4IWErc5Bnsf6NH+CgmLOnsYF9tWULX
Xd39EzP5kNu7VTxR2JDluuy3tnmfI2wksVt/4gx/aeudhJHLQlk/fp2Q9GcsccLxunr3bGSusJex
vVrd5DIaqiEtrEARBW5VIq6KSMbuDgcxEowTe0Gl/ONfj26wzTUMH6pCGQeQc+W6PWUhsxwkTSBu
Lpa36ZVhywzvwPA52jjoFsnQyWZj6xgrTVwr9jji63gZitg0ayuv43PVB/6EMpCHDVVzS+RbvAsc
bBZz2lsi8hBN5j725An1LLtEM1XP4pE04KSRY76wr0hUce4+uyHvlOuKjhr85V613fNiTzGKFML4
nfl7A7LFxZOomC0u1XXWIdAvL0LLNulMKz6M4iVJykacg3EnaZd8lIOFzfbKGk6daNyap7YxuVeK
viOJvqjQl9WZr8sc3Rhp81Bd334xTCX86oKJsEBdHQ3vX7JY+EdgpFithBj5t06ZCCeeNhLe+RyU
bupdDdU3iM08pNpFgGyOkhrRkq4HcJXFcuS7tHwp+xwmPCYwU4Y9kX1Nkxcwm0biZ+I9TnoftckD
AQv8tfypxqgzkK/sljXu2Y6FptqME9L0SpOFYTwILEXCpTYx+7wT8IfTMGMdNZTWLMHTaFQEc2yZ
Vvddrnm5YFM9f410g12CeoxUHIvghBKGBIkQQvMUAjWIS73Ak9waNkUBRK7B3M7YUOI4C0j4QALz
wx82zuaisuFNsuc2eEtxKm8hiExb/KJrwuvGTzaCchkUGHW7iQFKN0zA+0D+TceTsYfnyWzWrd2u
OEDY4mGa18Oy+4bnayFRgnfJ8VhOGUc+WB2cfbUT3g0XAB/UWgPM53sDjKrdXM01ZLlVXTzXUTxM
FJBSS5ht/ugHglnGT074VzKLElcaO4m49flB9AnudEaB7Ps7vLBDIN0a/I5hCqaT/RhBnxvP51li
+GA14qEJk+u3WOueQk8sSEcc9zK1W1WFE9b12d4Wo4DwWS2lqjNna1wY03YPIvdaEIkPL5ketScr
cijPsSVUZoAIospljQ/rfAFHkY0+x6008dALLDkcltfANocIOHnf2AKxzWLM/H8SuP4izMois4FO
NmVJf91oJWsDjwl4ZBrYfYbGOgMiWTFeEtfJDOaKDl/WIJGxTyp4FpCpXJSgCvZPwiPjNpq+S+Zz
sC1vjzPhF+Gy7xJWHAW5GHvRdzPYdk/enZG/iCMAaE8W3O0JE53S+lzVDANbP/cK+wq7uFPbbMLj
p8uLge2cAyGpJWovDxhK4ChOlsrRKxJ81dAH/5J7d8tJYdbjMwRHgGfpqfUnBEau1d57qOKUJuWL
v5Aw4H7hmGPRxRYNBkcreR9WotdK3JPrbJn7fmODqln2Nr0Sg3Lhmo+xTK9kMu/KOdpIY5EFyd52
hMx+w6HrWC1mfHIGkmYABAHvViz9KFwrOQKWO/NxjO+fNhWlrG8lKLtmOVjL+X4iDP1vgwwNmPHO
a8ve1f8q+qJxXgk3TQC4X6vOPdcS2gfb4RxPMZ0lcfJuCgT483O+isrHHKX9gzNzN9JVEy9HNOG2
rt/KTmpqVOt3azEbeLJv/rXm0HToyDqQRcRAcsW3tgk2aeJBLcuykR/RzYqDhmzUcsoxkcBjLjSG
hutiUfMjJm1vtsLUUPkcWA6eoEZf/JBwTX8sAcQOH8QCo7X0kUFDVUautqBSC6apGo3WiZ9YONJj
VlFvZlxMRvEy6TxX1stfuEq8xjrCKslVmHa1Oyc+k5H1VoZnrj5gN+ZhQfj9ZLREUJUNfCDQ0Jl0
qc0qwCOOxrU/s4dyV9+c2Emk/I2uxtvkeVaHzPEvT+bQS3SqO3h+D73N3nm1gC03aoPPily19PZk
lR5lVekbes0jWl9ZjQxE2pOgH54LlM1w2wy6G5hE9YzRgcUqBXDXo6zYjS/c7vagBe8Ca9MiNakk
IWzBLFFpZjCccumG0emoou+FpkRkdd8za0aiUC2RD1PGxh0Vn8AMXlX+qJk+sbhc4JJgWdF3l2Ap
pSNBlPB8bWaP/cr1mhXr3xPAKXUWCvuSjKHmQnbWjbYoQMZxfR2hz83eWwJ+ubsQ/u2MeOp7/p6N
lB+5vNRvLnn5V9EvBqB/QP2qeJN0cMuvtX/wY/v4D/Q5L/ZlC5bD0ykB9TMFQ3+4cfvRmnwks/xf
2R2rcdFAIacDDmSv5KkGVdfQiAtKQXUY3+VCINQp0YUGjzNZ7kQzgjL6+Y8Jov0Jvx42EkliqAu2
Ye8uBh852a0Wt1ag3OvnDs2rmx34OYDDFnJteeHvQFkxkZYRerjHkmKcpi4HnT1TnG9wZJqesUuM
sGgA2/UL0kqV6R8uAKBDCV8cZl4q91B5KpxgeBxLqVPG/i9CGNsTgct+4/jMuO8CRwYHwLm/B8aq
aO2hifY9dM7TT2NWwdn0zFuw+aG1PpB+NaPbGi3T+K0WypZdNGLwWC+k0/VSPhOxxtXYp/tOHRZ/
qd0I52DLHG2nfOf1o09nwTnrJU3yZI0TdseNgx6XomB69bTIQqEPEHp438kizEwjbzv61lNBSNXf
MO/4RWJzZHJ3yullvtbnpEMIPxdM4ZnnYkdqCyxa0hQkUX3X/NjjqAafiuCjw9zoMhwKpoUrRZNp
5HOeSsp/Z0WgzwgnO6opydYT7RMNs17Bu5lBGzljlCj3+7vI62Lilj/mgBmU+7klVTR9DGtqaeJ2
PnVrnxAgTxQsWRYAh2X8BslexxTeloxaT7VlDhTXe5Wx1ImwSn+6cxJdEzNR5NmQoiKmi8PgGjTT
Su5l1YrysV2Kk/7QSaHaZ23nmO5M8XAl7fBksq9d6wAUdaUE5MNOv1bq6smPgHln0LxdGVe6AIwb
GNne8PplP7sV+725bPT+05DVpytppIRiTrUtX3gZviY55jSeWUykNWtSgDJ5GASoCZitpkeSrqeV
fhRWKqqMt8rJsag073AvDkP8JQV6wn9eN+aj/z0TUvNvZKozDu/3cJ+RpFQE3s0KgwHdaFTVKA4Y
Lfl/VUhjj2JIedDxG41mBIvubJ7XjxZHIU0hxcAX23lfk/mLPNFY2UwuZ+o7katBQjSMnbYkd+YR
gmYyxjK5l0g/RAFlZGYtKVQloRemBJO3svYjPzm4tS9tBlbA6X0Rcgrr23TCoMBKSeFL1MZ4FmIq
vws2ezqzHBRhlTyIzwZIUdfB2GzLPEnLhfpNiOpPyaH24EFrP3QaalCcGAkrYBneN51siE2mEuNu
V/MqnGUzA908GdaXtMY2yAobirPcszAa4A79KfQ5jZLm6jkscAVzC9JtseveP+9UHkbbwZCZwnWd
HwhxqAn+atvNPaSWyPK4Dno6pHV1VQc0KUGGBdiruItZlHACUxkLRRwlhlvWdZqw2TYu/6RLYr45
IfkU5xgYhAFPHr16KfFsFh0sIFTPFw+d0258qfvrNerqyqmImgFqU/Gw5iCKi5lu+WEMXqPpNawn
WC1ZjsfaWfULpMxfh/5w5LvD00ie21RO7SNUJh7H5YsIBvfxyz7ZEspmV6Z/uxvd0lmEWm7tw617
uGWaHYpS7VZX0JWaH9eyHFyFut74XwSTA3MRt1Y3vCbPM0qDJIz0p30KKloCkNOSLk1BBGsqekTl
YbzbXvUFHMfPio7wN0HoOuWcFbsBZQbY5OeejwoYr8avnNCppi64x7RvHzfT8aC8qVhjutSTwQwo
U0sc6GwCvD+7jFYVsnT5i9Zl4F5Vb3f/OKFFSmpagPQ4V8yZiHWMQ2b3Ro1HbGPYQUF/Jbfg+1+B
KwYmjhSmsG/bkKvbOJnSvE7xtxnvL595MqJD1hsTrMZKTeJ+xYWM5g+BGIg38NpfZu72/aOoGhUC
1ig2C1VRFgX1YUUgor/VY70gPjrPe0laErON54/87G76WQ+l7Ps2bI5Tq/67Inu5EH17UTCwzi6F
E6xonFwDSorR6Voi5i9UqWvAHTyfYrTByIMnawik/ZD/cELOWHooP4EbsjxrnDsaOtpL8NDfj/LP
1f/tM59AHOs6MVcOscd2FpRAC3cd8jmJcgOnn29MNyy3fd5AGSX1dcS9Gls5c7y6da4xnJPHjWvX
a1OeVs30sCuHlok5HQJej96fQdNDoQYEYKwAXpnkaOGVQ5MA28mQtyiC4AZEaqhrY77bEfMZJhy1
9HqnOQ+wKd3yAwrcmIkRSUF/0Lm7M7JE+S9LNGQnyepr97sjbHIb0XgA+daSZZtVcrdUYbN7j/HS
CoNzJSjxNMwee3+oJ6vVowcMtAzboR75EVsVRM1dErD9k4LgqOy9eRw13SuooW+zGElTgvxRpRIU
T08LcnBZ0P862JXTbctf9jQXYm2dA5fWT/C3M0SlV0dMqdTdxe27qsWXy84eY6Np994EMiYZIK11
gGwTL+k6UfMVHgakRPX1JJ4ZH5cTmNaXhd/O7P5bmJF9qxGZR4VwsRUIgj8reZ0I9q+oJIPuveX1
Ggd5U45YF5ohCgA+Cyts5jREmUZE4OSjqhZ9FukYewmxoeLBnsD9bGzvHeeoIagV59ecTmdF7LPg
gcqKMSp/lAB/JuxxfcLMVjMLPF4EQVMGFSco9WFM1OG+8/77tI1U/eVNh+1QOW3Wq28s90mpubwm
o4yvMO1u+gX+LZkjQpcER+SnVkD2gMRYgqJFQ9amipR5OWf/HcpTPlbcf8jT7Jf8Islva/TnU5fi
8Dj7YSvRHwDC3VAtqQsNW+IOMZFfxvIcNf7oTMp5Q1sht3nKO64bLU6X435X7oQK2WvmIXbw16Gi
ZSo8cn3IBnEqNnA7nxzLhvxNN6lYP5KzMtvkS+00JL/rYP0766hc6AtP8BWYuv0/LTGkSoQExlKx
Xr/+CV+vHftU7+pOKN8SEO03EPBkJPmGm94FmgMa2ZNlONkc0S3fVR50k9tc4DDI2p7fBGxwBDAF
Qnfo+qfmaJliSPUt0vFhGo3i1H7RI2LBaRgrIiwoLii/pGdl/rfNBOgSdxxUwvLemy/IZZ6tmV0y
nU0q50+UttfyCZiJgFaK9xLKql4PNIkiTR41wx/TlZidw3JCHZdfbVxMgHc0cExnxJ+BAcUP6thl
VsutN3PNeVvT1WZP7qLFQaFP4GDJoENHB2EbRBOnibXOzrH1CC4r70bl9T1kyZwTZ/Rv2A0zsHj9
ZnO7tHf0rk/7nGM6YJIIFFmXlzzTSbpi87MOZ2Lr2yhYZTO+xbu1nPh0RX/WvHbM+96XduDGKptY
8MqlzKNC0sGn2YNdZMeOmGKJ1vXdHGHz9ZsB6HKqSe5wfJuOtG/7TRHu4omoDPRch/oBVNIVGoyI
xnnSXDaXwSUiw8NVq9oKVOUweDoHieKRusJgBdEHfO78QS1ZBRRgJI7CIvcWfqIJa3pm+OHn/389
SBdtfzuA6bMnj6CHhdij2TRdqTaIpZ9XAmWZueKwl+eA/RZAL+IGuCI8qRTCFSH6drMe+doRGFnF
qQxZOQkxFCtS5I0H++s2qu9+9sLIXK+y5TNCwBTolba6o0UHAfiUbexxOjj9P0kI53LEtWSuwZUO
G7IuaA9v9dFUr+gnVgymnZWXPrVIVZ9Yr504S5eC0XpUOAv1ZPjcSgM/S33ysDNckn1uppBvWukk
6wZ0PVt7poJ1hMX10eiNbyIbliLtdDl01RaDrlDN+KuR0kfSmJY3DhAe5uinvTEcPd2ovFd6MRhE
NiYDFy8OAYmdCq46/fiQ7OQxwaQjqhB/K+vpaGFFYvHzUBITwvzlEc9xXmWH4tf5ddeK4qvXiRgW
nLQSO7Cftcl7wkdbnWsHY9VaiP5KyCHrNZMH/XpX6N0wwk5TmisT56VCM+JhgxPxQCNo0DeGeOJv
DZFJD/mBE/GvY1wPa77xTVsHwCkn94MkvPH4At3M3LYRynJoFro0TwR5wO2vvVrn5nGsDfKYg5YR
mzHfHDc4t/H1VFIPZ0AlvRcZ5qqlzFeKUxbSF3ynBHShheALTg9FY3JwvUDGPWoij/ADPM32xOSb
IUfZ5lWxG9PfJ9RNWhHh3Y1yTXI8A/6WD9hdBCJv8DBFh8mXH/WnasnNIwNQo5ufnIBcTCKnjsyl
41YMYijWfwI1tW88B720qtfQ9qfWsF9AtEepTwYw8UsMjFMcT+djCTLmiQmqwgIY8XbIxWJFItS/
kljffYFITcSj5a4bB3aGEF/Le1nA7vFoqvq5mJOYSup1KTU/AH7XaIvXIAk8QyeJ9QzheMV6e+iK
CqoDctRNpZONtJRKpq3Ew2IoFW7luwem3ryLZO+/XCNlCM+ZzFaodHyxzFy1Osf+lFeVuDlDgP78
9iwLrGEjiJfjTIx+TiB5p6YFCOhte6H3ME59/CXw4W4ZFsoDTzcYKPpn5WElRwewRCij+6lwQW9f
LlKfQwupDdOMLJG/BZIFFQU3XJpwy7U6e7dq4TpDhpGEkC0zOxXEOmD8YjFPctLpcaF1u5LipFJX
YawlAagrZzWVchiHFmSKT7s1DgpnrpzhEgQ1oKxkOvG9oA0qdzzgqg+3incqJ6pF6ScEgiTwkmn7
fwYYDfPCnRDRmOqtX7EZquclVHZ66Wv4l+MXskBHPIT2Qiyco7WzQ/4GWNvq8H9ezTtJuiWkb4uD
nAMKmI4y3chvXUJWo/LGEhl9h+Q4kUemAA4vVvC2utraRWJJk5qURVpn20Jy6OI0EV+Oizg36ULg
D242FfYIyDz8Fc4gqDMMBJGf15WiEM3EAQkrjXE5fh7sB5pyRJ4FwdJzCQ+j/c1KbFVulLSPDD/w
OrLITn+92k5vr0TDvDDCfhmiUCcPb6FgVN3Itc2nHil+QX5DgqPqpeYg06ObVRuR2unbA15WeVNU
uumcWpE3c+xwK0JU7goIUCOce5IDA+9O3q9FjFYw/YAzuecJYBn9Wg+Cye1AjQbuz8cmUFnSXU3s
LdG+x97QACDZ/Cv9aZqNnqqzn15KDfgMxi1IW5WiyUpCmmE8rmIK1NoYHJcQoHHuhVnlX9n8n7oq
ZH6q+U3ZobUv+pGySKv8Ga3AAzj6noWIRny4P97/XCtPKgcxZ85LMfOv8ztyUsOc6yCM18xTkm3j
kTlN3IPO6BOrDbMFFH/xxEm/GrRNU7Iz0ncMrJnN3XCl+FaHRe8kiCgvnQg9qQ7oQzBWT5g4XJAN
cD03E+jyOe6VPaGXeQccp2dNVYS4RD1KyVx4lNOaqcO02L2BndbFxFZiLwBd2y20mS5VMkF9tN+z
7t1uxBhIzj2t3dlYTu0wDsB0yMqm0fIjs/cbtWRXq51i2m2RDVtu+a5iid8UtPIT8Gqvtl0Ozqik
vUGl9fuEVggpnTtFCtP8Rw+uGRDYJvlOSHeV/OhXo5O8WFLP9b070rvGKVfI2R0JZ0GqSVaMqiOc
MyUZiKrEBXncxpBtBspN0vO1hkkraqO2Lc74gCVvm5wpWItgcf4Fbuib4icpoGP6GUKkr/TkCYPT
xSsha9EOy9h7N3O8dKCWJyT7Ncctuy/JwNvSUYzfVK+McN2uFoNPvKKyjLhWeB4HPqoRWs9ayfha
w9Uj5WF1N6KUhZAH9ckUEsSvTWMLI3s0sMoiO0GHO6ukUEQr9adnC0DQQvLcDjNlhS6jGIVd3fyz
EoppG9+K84kLrfqGuX88NtKl1+Q6UZqZYEnYS/983c14O7zxv6OJNyP8icrCQL5wOXwKGq0hgjTH
zKW+OctDopFsF7JL2iKfNFXuz94nWCgUQCPwaPavhq+pFW2GfZwmwILSGof7dkC20+W0SryY6SkS
l/fcbcdXvPeh7Ii5tvYghaNfUarbhrzyC+m+4I1cG4IFrbHFd9xLSr9BCIjlzLUNyQSZ8jlVmOXh
BZDL+LTmeMhu2CQiNCmMC/aVHq7qIdRK3XwlHJIS0yHweabA2K47fyqCyDGecJBPPqtyOURh9Am2
02/yzb06QcHAKExgzlRWpSfXueogNFvpNUxLOIXIiFer/a/iXIA1C28Of8xOKR632w3mnoV6bgvH
bFuGqqDgLA7i8NN44nfpq06XJV0Gc2f2tAu/Va2pMaMBk2+MEewyOkOoGBD3sDaMpjxdZbpAS+9E
34C4oqquRj5DDW4vCDtFTeNBAb1aXhWYyGyQXrL8FqQbFlBJO/N125909pUuQaKRH9c6dOd+QZT6
y2tPe1qq5FHMoOYM26bOlo3kOFHvbyBWYNGxdPWEgKjMtDRnfuorbfvUsBqOpL2H/u3And+5ohqU
D9euD7ersL51lWmn7JXamE5vPXWfaaAn4TAgzhbb9nu2/ruNOX3SqCtmJr9rf78QowoTVp9kvdZh
xqlqJv9D4ldZxQY4dXQFcWMXz9FUPEjwiy47xqIfRmBgxNd1g4fqqfKWS1joToSiabc2TQt/Xgay
+tRcjBl44bo87xG40LfPg5NfyUQFoe8aAhmHxF0HSnwf/QgSfTrsaDNAf5I8QAu4tGC/uQqIjZ1x
Mx3xPvlF70nPC67N2OyW3d5bK5eGMrq3n2d4ZQfaxJfOT9KKLgJjYOxGVTSIb1zg7tyzazFMzMFz
7Zjqd9zdlnb1ASX8qhc1zqbyiNXd1JWR4PhZPqHEXIA2hms0gXlQjOS94BK4ViVrbIbdKTSkrgBh
ZDyfMKxhBwnUntyvT2+NeuC58BhDxvMJQxIPTiFdphCy+AcoGmptcoTV+5o0/B12aYv10kfTTT11
OD3uvcs4vbWg4gzRZT4s+FuQhkZBoHkQB0Kxt+/gPozE+F7eIgRyK0EkQfOZCdBZ0g/V933MwPhX
pP+Gw4iKolOAd3kxH+k/azw3fscwW2Y6pbY0UqE70wy8s7pL4bx4xjMVxC9m032QrCYPjt3Z+RNS
/0eXXbWPgsVFPBSgTE3yaUASl07zfNf7g2GDCIQOFoa1ppo/aFKKazNIIArERMwqwFjBu8kh4i5C
Y3DCz9OXGACQWo2em1g8dnO9UmHDZN0yGCUG9bGNiTpR4nlOhUtXgvc0GQGCFxS6V1F/WwFP4iK8
6eVBiC7T0y9VccmOjXIySTvW4uwmFrGPevylwNhTyBml47Q+Gc5GetaChjkNV913lxHhaVwfhf94
PIVV+5WctnTCEb8Fum2rgAi8PMe2u9kQ9AfB7CKCg6mXnf8dDIfFIC+apEASq6nQ1cdyegVCujRk
pV8jTO9zhIUMhPXwcjtAWwn1oJydtQUPtRqSvVp8GuBGvX3Cy54vodX23/Ku/fHWSdI04V6fLg/F
7o6zLxblhFdFKqqx1xJOzifaPjPpe/n2AtyF9QjMGSX9220HKWxnd6sFIdaYtOMtVhcihZu3EDss
D9nxC9NxoVFd8wzD1b3+z32RgSWKRVr3Lt28xTs+QW4SA38rJrg9iXZemWu334jvcmFSdlJvjMLM
ehg9jrXlQc+06yDl5z/Hd0SmYUEr3u6+8msJ7g0+mfXBRuomZJWh/oqIuNbMGiCxtqQGzCIeVAL4
rlGX2zhYw/6i5stn6+jxVWkB3QwWfiYo5D94hBxW8vYGQFnszD0/3Vm7miODo0pX+7d+GtvIidTu
j42vtCPx9zim9ys5JenpVU+CmVSp+58VJuTotddL4n3WmZEWAwBtjhIUrg9S0HWwY5bai/wto7eN
glAWCNYRUWXUr0+R6+zVjdTWqLgA+YfmfL/uYCeA9GFYO5W6HZ1JnaxfMLHJ7ocqaP5Ov3txEU0x
aJWozRqt6rIMDsMpX3RmeVSkNtHY1PPViX43QNBRhFyMbcnxLiQieceucxohBgxxNz+jOe8XmO1J
gUubHlPnxIiWieJAiL7mLt1JLu3GxEbM3viwE3PdLf0kv9rIHml9nM1eeOAiDYwZEQdTov1tgVn3
KEPmkqglv7P/1xj4gv9elK5FE/J9UBJR9qs9GSnZQSCJOhNujnTggbqaWM6Cztr+T7EIsjdAay88
GIXGcrUhiTd9YFDpCDWCB4GJYb/cWBHrBy7c861hJR1bcZhu96D/VzQxuvRJcLJkHGUHMSq2Sb25
25DAsW5GpFPVS4ERroSZ0lDbFJgZIrpLuMrdYpAErVWW/UTMziqw+rDLRbRvi2VpaPf2ssbzj7E0
HVohWPkJwmtnZ6u97fsTTO8VTIo32WLLN84GObVa1V+Td2phcesSTLS5b8APlydSW5NL5aqX0yTY
J0H/D5zLIdQAS6oZEM1z0f/nDUu9t6k7/0Jm7nnG3FeIkJu/Ku7Tz3lB1SjHOnry+M3vx/Z9P+ao
taNuU3RFHSY8FNCPTJby7wMfd70Xygyq1HK49mGQv7MM3+uySsj4c+0cWaHbkwl4HHL7C6X8A6o2
L4FcGgLAnLVkOmjAHoCv+g7tLF5aJmftHWj/ReazusQmpzW3/Y1Qgas2MtQOFEghcKb1ocRNqHZs
7iM+vGCRJT9oQskcbv6iPVJyeSJx1r+LAk2m8EclHP1LHRWUUzOtp6odmF9WPsB3wjFvxMLxpkA9
c5FArrQ8OAIoQR3ElgA6MKLu3zHU+/zXSvybWSFtbsKx8k7RPFcjcFyrvFIzBCG4bvlggelcZkC3
/pci4VTYu5AutAn8Jy7KsUmj0NEXpI2RsPCVSDmtI4o6nxg6FY1S8V/wVfs9dybTRf82LpLWmPZm
R+q2KXIJnX96ebkRonwfACmE/Hu+b+MRRW/u/NpEzxbzsFAxxjUxMU+RU7ekneYWtLsdQlAoMuaS
Ey3Ib9FKf3F7AOMbomOOuvIObcNYmJhefjf3I8gUp3DJIPqRIPWYt2O4/vr6CYg3ngIh8Z8FlTpc
jgNtM+att76WiItcpX47vWRgNlbYxDzYX9/XAUI3h5OyoBZFpp9DqCbm461ZN1ZUXG2S2mncXgdz
KIimMB8swDh68GVdlVUPAR7rS5Mn8bVM+hej4DdfXjsW8ySsldcLY2T3kw2G1CwFgDIqb5mxb97u
Dr6DNfamtbfiY69bU2AX+Yu217M6vYW/ucfUKj7dGBb2pac+ePodpF0LYTBlGWlC7ILcGdxF6Td5
LM1L+pbePbURrjCOiv1vth416e6O6kETAilS8OLrY2lu2/ZzG86JNypZb5qiXNoB4RWE3uAqgxO5
9OKtEmLRpi4AaJsDnJKMf9GXEf3Eol5GGJkuF76mzycASQlR9J2/hBRrE+UHNgnras7UR3dleZk+
t3ZFEZ/Q1jpNwJpJYjHsciDtaiit+AC2KcHPEQ6I0AP/VvfQV7uAYzVM9+fLuCvoxBwVeHPJFCXx
Guv/yDseOExSLdcU6Zh6lYiaQyPlNma9qwOHNYiKF/hORCz2G8Pc1PflTfZKVzf3wPKAcNcwotbc
lGeKiJAauuo5ggzhexJfOqsC+slEl5Np8tu/o8ZkgViZ67B4R6G1kbNmp/r9tdvfuUcAZmHt52H2
DX7woKL+yXVg/UY8l00Snyktc/Fv8TuZ6Vfur7TCWG5OZ4gn2z+rkyPEvWrHee/f9jIkTYMT3tQP
+yjuIP8NP33983SZ6YKxrH1Hr1XRNNKWbSQFUyaAv7zFdYm/xfZKIoqLi7khE/NmsGnoHY0v/v9y
OtpAHbVTZ8rBtEVsIN6P22/cfnk08CWX8bgj+da1vSxyqtfXKV3YS29i4KSeVbb3e8lfu1DhBFSb
mNaxoV/nAnhNV6LhQ8olSiDZMqt+7MvkPacsPaFIp+KX80U4Vgxa9qVdV1lRHiljto3aIYywhEi/
h8hH582euJpphOUdd0Fo40//NIXCnrq2PkXL5l5pnomTNAdxrnrJ6PGz9K8R1dbW5bxn6v0iMGeZ
ifI3cNhcRfd2e7VpSDBuMM12+DnkZ1dMIjzRzpC7u8HeYoa6lff0+/2hJUzGnhR/sII23cKWHKUF
FWSolGUI+wVOCM6TrPIVtcu50qSGI0DzI+WxcDObaXvxCLSz2a7iPnyBVTIT1MwlBwutI01mazP7
oAuvFNuNgzdkolHN0Zrgcg5tD7qArAcOdhyxYq58FLgvXJmoB5WYLQ1v0vCEoHZsTfDrtEPhBbM5
clN7iEZNGKKCe4CFxruZA/jf+hz6ArAc7ILncGlgg6YdZtdJRVOUPbyU5uC84UClEu5sikWDCfWw
URb9VKagvfTW+40PEblOcqzpM/Rm933pikH+W6nZFQFmI54JCUi7jRVTuoIrqgslVI5KDJyrDfBz
ypSGphLd1UorR58KMY3WmYdgfJKiBu4ATnvuJwo5SO0V3ZlAG6Pr8yVbC5FnDqyaWwqDvFL8u/q9
Qi1n5onfYmtI99IOCQpcHrVKGsABnsRGLO7tROZYBTBzICmTT1rav9MXOZPRA8k1uEoWQTm88nyd
4vDBzjiNez/SqC41l8ewiFkJFzVZnh5f+GFyIyJ+7bHaPYVvvYXffKMeZV8vb+iWm2y8Cg5SjUTx
lKVe1juyymDUU4VIYLV8DKdXc7FJaGSnLHqL2yInL1c6QShhEBasxQa4ZEOUX9Be4Lz6VVpr7r5Z
ynyvqHUiAXYHEEaV3c6DizABvWNxeKbjg/fGwCcDVhHzYTOcBRIZFIlXK0yuTg+53I/T+KCR9Vaq
a9Cp0ZyzIjmQGlQgeR4bU1C3JwPaaX3am8wZeVG9uzh43Mfv0hRTM7NGaPjf/UCP92ijzFNQeV3O
TOOFqAd0x7DHgNUypuKr+/S7FwGXQFrtxk//WDEBxJHViXa2+AtzCWg1fldJg6+gFzBizujplYkR
UC3GIHlB5aj0+cnCudcgn3GueaxMoiwMXY8iOBvVq3LWzFJR/VxmIotBBwFJBh/87Uqu+HjfMxnj
8UeEkgfNeEGWGO/1yXy1rJgAYgtW6eQjce9f2NinRxPV7LC6E/Jb0JkI4Da36Gky5KOQX1WFndd3
5keK/KgeUE3KdPkSEYssdbqyTgQB7tfVLq8subMh6gXXqehQ3Bckp2DnbpoiLRSDeqC8zyKRPdxP
h63uAW1Henf/ueKRu7bxejQOKinK5AmPolSX27xJUQ5etICsqgYGSFl/+z9XT5duxFpGDlHGw/GC
2RLQPrfjDD4rrlNgRV/86vMFSmJyeTMb9aRbY5avk+kCSUZL+NSwHKLmQqVpmu7ewNa3rWv/FUl8
xnYPZXTPR0QaytqG3vh1JzT+eA0cwJP4eTC+a0QhQrGBgpYFo6COgDLdYSP5ITrGl5sL0z7hCS+x
qTZdplmbZUwnUK8DtfJBcom1yomd96guz0g6oTGN25XYG//qovNaZ1c+kVHzoMfCzdoCJFLR5NDT
ljy7Z2e1egtDBoPpUENkQFPSY4SBL/zSBmyV8MljKuUPZa2lrKRGlfkWl6be3iyjW/0Hd71ZAJSP
yV/wOgqzprQzTW3ViAvjy6a7mAUN3PejfGDCxB4XuNldYI3zJvHjZwzxaOHvaUFQzCZfz/8VvtZD
INMyzz0ppicWU2ARw81p0q8NpJwTRuktsxrEI2wg/Il9QeeAyPm/Tes5S+7EwOwj6UIRF1XE0hZ9
+ClIePhWsQZQdhI4msu9so0ACkCyUq9bCWIaJt/k4iTjVnx+6YiWrg2WgIEyueLuuj7u8X0UUwQh
uUeWrP8xBlXWfljzOAm8VYEPQfGAPr3N6bim0PPFypo+fObv7UZHOTHGox23YnjOY6G4DiZpPaYC
Z7/VUq6mSBP0PajZZ4fsmBCdbvLL4vCxBJ5+ik9UOKtKB09z3IUoAOtxboZKUhjnrpvrAlHQDBLm
IrvaaEihLFhujQGdiEyZ+fuqCL2iYJJgRCSXwXHjLEXP2Zsq0YYKH2TKNQn0xVUEM6X/INLjMPZK
zCOSgc3FGDoN/3sj9QfzjMz+JKH/XiukmTbsSi8PL53LEq0RNoCBzQqJOj3jPr7t0TUQSqdKuEr7
kH1DJA1sdBL+1KC2Xr4nvVbDCxjnwcuMp/9G8d9WZKPVKUrAktvUQ2+t+ix/2w+ZuXTDufqRdfw6
xkf7VFahFd2f5JLp5RdRU7/7RHae8uwgEFpz/x51Gy68EJQHm6RC1pY8Xdu406MhOjEU5Nzpz/LV
RdLVtykPYDJRdG8rQZjyj6qPghskHWF1OgoW6GrvH16XM87GhGxJfvDjn8emdbCrC0Ay+AmwLCfE
2/+i9X6K2bZsZEaj2fVPXyMc3bPSthfJFlGcAbn/0KKAyeZGmH290cHjIQHtcxyjNPR48mqtAZlw
xDveQKfqyZGdQCIaisSzQ8X+9mFwXLDQCYXPn1Adg623yNNziB2fK+ulz1d3f1dctxjrnxGGuy3a
H7vZKmsNYvsH5pWSuukDkiKlvoy9lfcWLF5Y8PwqP0YVxQzgCpb9EM5fEKpeTgBM/jGzUHD+3135
9RBuGDiWDQXmCXhn63u6IOIKyTD7j6/Hc1BAHvDTV5xucRsoGkgWjfD1fxuqr4nDCas8g+cBotun
8qT1O7btW3PF1jGCztUq4fJfCKElAUuh3goVgiONOrzh/Tb/VIwlm/m95QhqcqnUJ6Ks/pq6MtgJ
JpShjXxmgi+wHhYZBWb1MxHkLHdyIkTK/DAyEweBWzltjs7EnpVUPcsPkZDN83MiLnBvMSHEujT2
gbvHGoAKOUOO3PsAQfiYM3PzM+lsn+DAn3wu/dZz5VNJUYKrWdZcZxczbOY7qxTFIN7BJLJc+QUp
yD322jcHW8hQp0Y2HqEKjC6wzJrRSFr5H9GPUL7ZAeU+/+XLPtNEVsylGT/WCue1gxPUZr6SSwPN
muVpX+IsXsRTVe/fC7iI+mQBGeWft8F5QySzObGoFg7s9ZXzvRs56QOxg9LZydghT3kVEZEPZk6J
p4l4GEUTEh9KkU2ic6hjmjYwBFRUCFxasHAtyTZ68D4nsqL3NOLvh3Rr4S5glk8SZLhSrsnlpsOc
eFXKdxuqAX4hm0+JNB6J3NXj4VHu2PaWZp8P1MefWBpIijGhyF6XmRcUadTh2uAP0+hVkJWWEbTO
+kLVkJOA+hfo2akqXh/M1MR0rWQ3+pW7tgOoDg1quAIKvNoRs2K1rK7kKdXF91jfDuzNw4FgRvCY
nrHubLLOzGhSFVQIMBnjjhfUejh3TH1+iYtxzFBwHdgHw8yojDxxRBcojeZB8s0lvCvqekv+xbgq
ThJ7DpistOdCNc7yKLm2ILOI67gCClRd3MkKQ4kYO+5kLW544i6Ao7DyFVdaTLyHq7TeM45mMWlE
PJRuoa7FCwPnTO43BmdNihzHDGSPUHO8X+Jz881sD6RJ7jKDyTMH4QCUCumVFg24xvCUP9W3IPqD
049+dvjEavN904M9EStn3mMWnGE80s5f+H2V2kGxUoCrfn2N17MMzD7L+9ouTkebfzeOJo12jLXi
XfJWFlAvh7tiEZmeXYNI+pua+lyJaMNRH9GvxWn31uwWNgQgaofIkzvQByscOv0cvkZqXsILhFo6
8cfoEcsUxyW/SD9LVTp/apfedlD+vNC+cfdqI6z34WwTF8bAcdfLh4o0nAIv1QwAmokwCliyC7YF
Irar0r0yAOKlBb9RSYtLj4hJ9b+/Eq5nwZubOJc2mU/CZFnvDv95O7v1QGZTeKDBnqs/LGSr+TkQ
bo/SOB9UuO6G3juTib//PUZwfaEYkmKASyMAdiKH4qnCxrnOd99GlLX43TxuCcNRY1LFubXSn5kG
nOodIcGdosusswmqzti0lnpCz0aEs9UBaz8uE2esWVPNC6479BPks/Ks1neyB2uehyUZOEp4xm25
sZoVtLlrh0JlcwU1NUqVS7IXc+Aq129Vreeu3lMhvju9CIgZSh3hd7irfF4ToTLE8IIS3QJrw3lS
hFZj2m6pcm/4bnZdL8qwSycZULu8MvnLAbSfmLC/B3+nol/o99nDRwvmvu4085jdDyI3Nb2nqPFD
KHDbTKRVtqv8mtkNqDH5AGgG7H4tvwZWucFE7WsTEa1nuAKLdiPL/F4inLhl9ayg+quOfVca2tds
e0KtG3coZcAHkqhwXg9aZjGBPJDGQf4kBphhgx39s+NsEYoIvfftAYfqPJEq9sAiFeiBZUAEqoXU
WMedwIdOuzYBmQA9biTjP+415GnwoV3Vw7yPeTwCbaXVjAGr/+kptWgtylBFLykChj13/WyUP0sz
3R7RL8UTqhSlOvS6p7eD+s8DtU5qejO/eYuSGZdu8X0+DT8n5npLujyhehn1BMlBu224XUpBaUk8
Rhw3tOw5qf5fD6C99N2yGtewhZaAR+mM9yzA2FAZ2jWH/5eLzC7hDHwSaD12zKiTGvoJnwl3g5y4
m27LQz8EoxxkoRlkkenPQZnnAmKgZOOPr8dZyWq5b1KWTeZpTvct4y2pnRbrf2aMR1c+nXc9ENXD
JVxHbRqQO7PcXbfwHwE9JEy1hgcypRUmJxPP2oLpzs5iXPPgt6Dgj2L6RsIn1iJdarpmKYFH4lju
Q5UQ4jA/8/2B1DVvCcJlvAiNkELQWSiDBu+464o/i8Ngn6H8ntTNlyYyks07QaxnOOuqJl4/QQ2y
z+r1bdV0yv1QXPrxrxysXpHiadrJrqHffjOemVSHfQTWx/ghFcqBCXZOBHoSqFj75FTuX4rsqze0
NwMjJKtw14C7XRGFkkFWqZFnGmDN4tWI7Hx/64jHN7L45Qz5c8M+4VvTH6MRy6T0SKiPMXIlToCL
uqvbfghuXsSf8jiDQaWJUYTmMkTUqNmVFq+k6Er6uMQHDSZca2For/1wLxE2DBjHyQDP34S/4xUh
l8e5oeFqwj3IcfYE9cMlw6l2pIc/cnvzY1k554PnzW4MumAU5dt4qw0RWYJ/VoVaBCTVXNCXiwO6
nHmx7Q1rmVLj/0Ij5X5hStCWQSQRPriYlvALEtmb7KCDArtEtJrBH+ix0zLNDalqG5bUmpF5o0bD
Mx85fEi952UtJ8c4PN79rMar1P68Xf1AJcYEvNjKZ+BDXhvS9MwFzGzIURf5ZKroX+l66AoEpr+q
v5afvy+9bDE7Dr2MngMW2vKCLMSJtYtBfXEcd17z0MMUTTdRl5AX2IR+aTK3taALRdZWSxtFxdiw
LBtEOxlEis1l0UYdp1jhKyuxBeZZDt2pHFjc+nElj1oBA/NI6PjEL6WU7G9KInTpNkEwNW3qxOet
jamoCd4Cd64ydwUwm5uHEu1KIo8A2uKYcfRgK1EE2uh2KpWF35TldE5kHLsu4xbe2DdZlutup2mA
it1AnCvVtRcU4D32aMKt8mCDTZ1aNR0Jvvadoo5Zo6vembZup8WuXkoSoESCXz9Cxqv4XMkji1HL
b7kPxD0jthTzbaACFBnmMFLzjLVlPYI/K1Ps+BxDl1V1RPtWRMjmmvENMKO24km7p6unye9JEfD/
AypTU5sA3lC9cFyrPEqb/MLj2YTCMAlRvSShMeQ5W+4JJ+SKjsPv5md5tbUdCT/7WQSWlYCmkUfC
ciHg6YFm+fKuY/DJ/bmiYRdE6ZLQFYjR2HDEdNs7HUiWnpQgXjNhuNi+sik+8c2o9l3PnRfkrVhk
ENn8TcXqI5aWUOBi5yPy25srxUup7bk5ddys2hghTVyFfXueMYAWSxj0tZhGkTpQtOtsn4jQ2i0u
uMrDxd9IAHktVzs1ulWEXGdvFsJNl/SL152OqsIBaiCSIt2DeV6f58v8l0QT/fARHhkxfUOY1rr9
W91Wku2/gAZuUfiOWVaxC28z48gj8gKDrouAkf+eErYD9Sw0Q1epiSnLAWFN056xjsaLSyMUP7hp
+c7Ahm00gNiaxq9cDKOu0e54CThbu/ovoSA2X6qSKLZSRx3w6S7jF6cnsguOpzQIrIsLcO2MVw8q
DEVCmDPn26oW4Xxq4Aiq+BQf0h2/srPPhP+/TgQgm1/JhspkwJ5m3wA+R7eRFjYw3vMeMloIl1qk
AE+vrbtOlJAPrWH/iJxKBgZiZMfyZDozxoZl/vJe6qf5eJqQyyiZS0wa+nzpBW45nGSYTBJ2wtRw
iZWRLQ4Knx26KSctBQMfSbrn71PfM2zev+AsqhhQqksUHtE7eksxU169y85jrpo0oglMt80bU4C2
DGMybgiSm3y8eA+glw/loRyKVqIHDdELdkuI9s9Z86ib+w9ygye+8L8ap2qz2F7VDdsFh1+2I7Ft
fHGoWt5blTR1ZVB+HNbnkGCXrXFsMVIn/37H/yCplbH2pN+BlaOoiql3LhgrRnnSYnopPTkywF4m
jNq5xpKih5OlUJQ8Yih6BqGLuLZgILiNqGs0YPPvnNzFTLS4f8+fcq9fYINn1WKMwXb8Nh6FRtFE
kEZT7GoPlqptDdy+4/fUf207gWleti1r9qvxB5Y5sDHz0IIY7qOn3LHXUXM3x1P6rUyjdI2mriNX
U0Nu0wXN6+5Gpj7HhFfPZMlOH1qVaMcgiF09fqVYsk63ODfA4bSyRY+trhEJ6S1yU3DRXzPwHXzg
Cf2FBkB4/wziIc2No96TIVgVl8b2KuNay6uVwS/64p2QSeSEi4LUJQNYKdZz3FCZIZNaUtATOgwl
L9WVYNeNWqkU3HhBAMYP7jTVxtBgILj6kDDjgat/RjA735WORHBepNTlOQl10LHiMbez5cuOFF5z
Q1gox4It7zOzKOtYS2QtcFZ6L60HSiUfKlZLl2fA+n2A3EoPgHNqTf4UnvcLTY3cAkuGuzKD91yG
3xKicPP2RPBdGLMWufkOR6qsCn+BivbanVyAjx+g88DfWGPC3E22WSKCY5YV+3H5GqGeNe4tryov
aYGOaQENkuCRBfupp8YKPd0ivL+RRNe1kgvgvnDSqBa4xG9EJDYxbZAu81OG7EH3UpIgeJY6ilAC
08B8R0ozq+VUw3DkYIbE84ETT0wKfCSObbIYtSMgvGO89oXslLSMa6EOwPQ9GLDjeeDQTWr54wGk
P4+Mu14rUom4m9FS8VFCaksdoanfzjMp/Lid+IWZnG5E4ZI745yaAtLA834K6txELmZc2bFWHZCu
iQ+C42578qTXZG5H6vyHDYBmKEE62DgrCEbonf4AJy8jzECyZzq0I+2ChwGAoQ7zQnpgHxA/P/QD
jcN4zYn+3QscfDij15Sir/mOjCXyMmHeYWWBLsjomuem6bncEkBBTJplNEaLtw+ag4sStHD0v8p/
nFOdksof/AFZuDGXk3AVHITCKonyToR/FbJJjnxHujHTg+ucp5hBoTzPeNnN4T23zVwvoYmt4iPG
9lDFFXD0JDHJJDP/hrNpwH3bC5GeUE1sH0gZJxWycILQ4mAXX9rvfkQPN3j61drRi3ynD3iTbQzu
gY0HcIaVPOL/2OhRjV7lxoRpo7q5dSYguK/Smg15K4gHKn/bJMwuAkVtQ86tQsq8YsiSSlmEeZlv
9yA762YCMBn2Z0mgsCJd7a0DrQ8rtH1kdCjFXmR2PQm13An+Wdpqoi26MQ+9Z4COOHQOF+SbEfpc
kLgYFRDpjIxG6XszcG5w/mCUV5L51uBI0rzAZVMokg5h+GWH0NG1IgWQv7+4U+f0oBmydzHrvTR9
HkMxNYSiJ0sM/ifG+yTzn4aB+3p3VArXE/os9chRqvGogMryRrVzAYfPPzq4RVSCaAiKVCeZUCTY
ES1evHNtYZTAIuqByjIIuk2nFhUdHsW///SMVc/0NYtt8Lj94TtzWwrKtlSYM+SMa1LbdTFAEf1O
IsM+f0v3NsGZIMqxWRAXLclSIWN80HmWBa1Z0Qm9YPJ7vIl6FwMRiRiKaVC4vlXOhelTv4hK8gVJ
5mz5CzIfptXKgGEPDrmOh0PbW+1AWwm+bTWZKSabnfq2+aLUSlq6tWqrpcNKAA8CA/GlFqJaUsQ4
r+2Rv+24sZOlksfiyKK4IQwH2KCie/AGGY88mAf4to9Nl929FDuJK6B2dDjFaQCYmtA/TjhdGhZL
xM8a8w4lpix+WvcsA7AJ2w4Nu0YoOra7e8ajE+sroHIp81Ju1T5aEsWYPyDmDkqWNqpBb+NFnKrT
jj4wb164+M563S5vPRT/Csy10/wW5KhI7Zz63YPU7QyRCv8tGU3uPf5R9SfEVHrhh0uxV+FTiiPA
ynJhzecy8on8WHQcWLnzWPbtoNbD2rTNEB02lTcZI9Tr4MJEKL82owSOVvlpveKk7yuzkhT6RXrM
//ziWquCohY1bv+TzkOHwUZqzWmgDAHH7kvfTCM2J4EPNDXjCbCSN3BYZnRx046lFI6X+iMET//b
ekquN1TscVA1gQBfE8ak7rNKfaSw3oCo2THPaW7YiGzQipRp8xBe6Ts4iVe6pQSZBo7HZlNsleJR
6lVHiCkXnq0RK1Cvxrgwlhxuvm4mDhDHRNfh8rEorrABpfb0CaiXR3+/eMv+vBstf4c+ov4PgfYj
Q8LU/6mNlPucrYOqAnr2DDFm7Ung9iN1RtHrQjiQF1rBNbQQpU7PASBd6FzxaqKr5pqZK+mm2HjJ
BgiRTFiJVV2XsOVF5znEcfC5C23QHwvjYuwJiwOlVXmruJulHA1msXlgQY/HNKXWgNNe7UDFZsgp
uIhAGtJj2L+p+tQ9w0Xin9vghdTKlPsXdTtODgN1+TaiRnkuQ0C1P1gzWOuDnIX5FmJ8BgihIrgt
eH15nHI+rejCmtFi7rCpDDG1qUhvf7moyfKbOYKSjeI5ENRyFdTHtBGjMFVVciMy8wDOjr+P1u8j
CJjbxh8WEtl0tUoMAKken27GGjCIbYQW5a08vEq4lTkddwGlmZiVJ1OSEHwGPEfwAz9GyZr/G1gH
rVKhqmAUa9bNZN1DtLu05jAnGc/9HIYffP97uYTeRvMj6GCIIrNmuRLArwZi/SQA/R4GO5y4SzH1
GWRWYkJKrFIGRkHuNXSWHel6an1Abaxdf3xt0SA0kmS16iGxdkP5xnHA95NR9g3HKCjtrNm04FKT
olauP0qZYzO4/ksNZsukZNj4H7APHLoB5PM218IyA6KmPlI2anNqzwseT6uiEk/Q9OcTyUzTb9+h
1Zqjob27W4eUjW8gJKQIC8PeoWLb0dA1Zt3AKQnHHOmmV+BYjp0TMcn6tbYWfbbtHUjMnBGXYcBB
pmeH7WS2b9U/M1uXY2LBYV3g8Zzi/UtaQrKYkoLnQuBBscablKgGdoxTwMVLv90kIp5yG6AzLY0v
CwQxIjPqEii0QxEUV4NLvQqljX1XfhadRS0ghKyDdBsFO2EKWF4qNllnm3uGu1zmnLsF2T6SYWUy
NXCZkhrzvfhDh1NOcVrppiIz0vrlwPnhM42Nkt1MUpSf8++UPmHbtBWuIxNuVUfk12o013QD8WhP
WgOVicjmhIjtsO6t+Wbe1vlu8qtraXfhRCoT3BbqYYmI4tcMhKZRhp7qg5qeueAB9mLKkZTWxm8c
rMAz/FPdvlQ2XL7s/uQbhdJ3/Cc4uNBNyH8wwGWOPvqN9A/gzoBPr9GeGDHUszwSZ3OOCldi81Ol
brVMJH2a8Em8SZsgQpVLBRlhNdLa/hLOIZPBbgXA3BDHCt/ApRCGALYMAsatePvvPuuy5YzSx9as
iuKbmmu83Wk9HYQOFvGoZNzlAXbrM8mQu+QUpmvKlZ+PAxm9JC88ZoxV4Sh2b4EnR+9xFeauF2c5
yl1YmqgsbLEWXn5XW9tJK6nAIiVu4Km12xfov0V7769RQTMdv4DOYabgQTP5NFvHkn7PTImAqinq
RM2ux2u7WDHTJnWW7dDwsgmzj6ymE3WIEi6PvOeCwG/Br6uGZLGR6dT/XgtmT5U+5I14kREdhR5T
jwvwBcPZ6tz8W8oIskHjQ9Zvo+Ve7v2KMaJTJ4Gf+BsH2XL7UW4P5IT7NWVkNKNHSBcIQKSD/kno
cnTnM+w+YQF8FgHIaOO1vwpIUz/sPd9cx59aP5I71v2oEHMfcDwUShr++VnpN0gY0LXoei4FfPnV
RcCn6qtRY4GCeGGZrgJF/ekVoQ3XAD6WgI57dWgBt06+4k9P8N6Zd8+SW2TsaqqXRucyMUOEiKJK
SzYFv2RZfiCYzYjAKwPvUD/YN0u1ygOZ9OAou+67NOLTLfllB2dpvCXR2UzQvHAIUupt79APV+Hd
ows6eXkLIK0o2iCRPPYHjYUAHBU3HNxI8VICPA2a0UELyU8a8Yop4iLz14Ndpflp39ekSvPTZEWc
Q3JsxzrIzi/WPhlNP6pythKrxP3HBtFOV/ddYtMzfFug2T5HSAkDzk17ZdMN2Llbllz0U/IKgYE6
+t0SdQHywhZVKjPyjq/35JYpuIy/YbUk15rpqwY6Yb7YISgswL3oz4mk+VrAb8HhLUwC+fTwwubI
gas4lVMP0Lr69zRwiNpuCny8sVxyW8sB95NqN8tSO2OKBfMY5j6yFYJcYkJam7xC5o25IOfIGBOF
+lLZ2XWB7Cl9QTbj3ZdBt5mmBl+PAI4H2F4GaeQIJT2AGkMiJ0qPgqzayLbtuGaU8oTuLXEKhwY8
HqnF1v7L1Khr4MzgHdLcNLb1uJu9phPYVjxfuEQlc+UvSfKim60uAgwUNCO+olX3AVyokpqTa3eJ
fOuoKBN0qBdb2mc6pKQWezkYAh/F0XHUc98YMHeaFSS5IZRegRqH9H+AqXbRkI3E3eMm1xpdHlz4
InmjqLaPEg6nApPWZ1WvWFSdiNdLg7IxsG6U/NDbfhO3ZSlI2qQ3u+dwAdAx3XmypsCESzXDd18r
nJpM0ineonC9a5QWAK28aMW2PyQ0rqwy8nSIL1C2+cdCiUovEtx8EYZAChdZYmrXiX5XhPErMclu
MD5bdzhLX1UeaLqF78D6fDkUMeDKF2N8+nUYm5GNf4aElHkRiF5L52trmMtsLWrN7nT/3ZqEj7KD
2LBwakDUmKdl1VHn1sNiJTa3Bs7elB6Ye2jAuWo4g9HrxHnLUhMpLOKaJWlyKoT9PyY3Uf7U8f04
aK9+F6viYCM6fKhqNZ5J/GY3m+Cf21GRRKpR16e/IPwG0UQ389kh3/kKzaM+N1KLk/qOqllhWUgL
Vu8LroX/ODhOn4DtXAd/CSCFBxS8rycMwIuX8MFSOTssaIdiZYVBD65mX74aekKFrkXHgWU5m9hv
GDmPJnyFp5/EmMvaLJNGqK+8xWjNA7uV10bRqrterP8oDOQZkhU8JfF5gmwD839ttLKctCCNrdGn
1x78DrZlsZqI0yQACVDmCSD5FXRWXmBtOborCzVj7Db3XpIlnW0r/0bZiWs/XI+9StT8JO24heW5
laTNqW0+B7bzfQ9liW3mAzMG6mCatO4IArCLFS6e1gia56TGBRPM+T+hLisj78jjC252dvNGjqel
GtlIoHUn7mHUrIediv1MY80dVd6hT6wGdEH35kz2w4wfYqLBgp/fhlhwh8X2F7nAC24GuFPCgr/g
TXUpFnUlVOaKbEdF9dtUpkVbV8oSmAa4cwEsWTHCHuB1d42c+oyhiBr7FKb5bnEgEMeyhOgNE4l2
UtBd4W9kgDQd73NNH74ghF1WwayoZq6DOhI+0AZfXADx8CylUQA8YENMDztrxmG94uIfdaBPnVY1
jwtLqpwi/VJRJAoOzn5/4TyMuzBOTAKJunmxR35WMsZr7IPEsCvptAL9zl/b92gLUJiWC3X/2xcd
fozgPcoZVfNmlVdGAVWy2HW7bv3RW0Mz6Uqemrr/9nF4xjsGE10AvXOnZA+aQX15j8faN2a5gJuX
CL4VNSiiFugADOirl15Lk5Z6XbB7kl8Mn9i2rjRHUJb/EDVZ53A/uaF35krJkuDQiSREEDpTtWOO
8NedpHsomgZopHg+1CkNWBwN8ZLFlSuTs0zYgjdjb3pzh2+j+LD2N2VvfPHhRI0H1JrVb9w3QKsQ
YQv1aG/F6Y1+mP2iImuZDG+elcjAxJTs21v8LqnakLi13ANvUtbT6S+8RSexdK/iOu5jfnIamMEy
a+s2Mihh14fON6PoAdXZCQhuRRoGxfx01rs1S+K/XcKjPhTyZLgGywLpn/g+S9eWhJ8TQRpiNFHX
F3tm31hmMEK/fIlcQTTbNWQJ5CIpKkF+htMIIh2Gs5lubfMV+MD+us3DrNvDVVjeTnnGYRTtxaHt
2GVbjNdUJY9XhXDo7QaTRTKyPDnpqx60mX+sXyX6HevuZGQMIULaIKEm5705EhFCDYWLMEC05NTP
IJJ6LK7Zr3j9NtYq1HPraByVoYKZkPfdYEbIBnIiqFDRWrs1w8eGzj8k8xcfA3O5o9c5jb0KIBqk
h6aEhFULcCMby7Jccx0XeJuFCnD6JD6X2YVR14tyr9uKC0gLoSVbCDgJlSkmpLKHWBFmJ9/j2SbI
bEGAAAMk7ElDuXrVHxEnVM7YN09YTpTmbKIosRENRyTQXu9XRewr9ZjYzHIwTER5DS7/q6u2ZixY
QrM7c3f2mPgoGYrWijiWXyyFd6w6GIH9KW4OGLABed1lbnQLc+/WgkokZy3LWeGNjEVPdcSyQnWi
jS96bLvni4WJMbzRW6XY6KnxfuFMdDpYUrehzbGRhi6GYoBH8LADOplZ079wfx0y8FucZAzsnT5l
X5UQMV5ieyK/20z8Zzlaao2fduULtgB8NJGWlonKwyOpAEGOKsJQtL1L9Wd/j+Sqw/CtPYTVr9Wq
uQOZLZuQqRyikkJ6DHTeZyOMovc4bRmMu1XGJ9eY/xb9UoGUsmUwSArB+XRErGoacaDKzWWIICIM
AULzEd9b9MEon/Ui1Gg9KY6P94yb6Po6vd9yuNP5tNEZ1lILKFDc9l29nkkMWmtKLffVPeUt+DGO
p5coCoLGpTrfhztDewq7yEiWiinv/6bHGHPbI0ZFg6bWYqJnMAJqRKOZtYyKD5W+CRE6APKhd+zB
d7+/bwG+0RAutLK79heh6f6ZpvKXOWe1mMo+IalCwswUdlpJwmVEP8PFa5He7x532zUL3+8n8vOQ
Au76wqUftCMOickZRJ+xu6EkggStYsdthScYCXsK/DfciG8/076FzTS768QE11oEc3ZHePs6Xb+R
OpISAs+OAhpX6a3tUVbjqJ0P5HFJjll9JMQ6ThP0UDliwKC+di54ppzRjsTcjI+I+6R/l/+rMc4R
hrb5VKVzf19vLcxuYJwHSqSWdJ76u6BbGviK5VzTCu57HYcXjq2AUyt74jCQednqaay0+MhXxj/e
PmtCgB4yx0psNxmJVxOO6Oepn1TPKMZLRmcbdDoypss3C3Ys7VsSjKXePdnZmAMRsuG8VvPjuFSu
ZBwWM5IWXUdw18PUeOOOg8/ZYHhz2uA8XfuhBZIS3vT+W7D/9gvus22MBuCYZkQsJI4T9swdpKgw
fhnaQYcC+2fg9CqnL8UDCU4dVynHNDfdSsBcw3YSH1KsNAlZKjCHL/XY8QJAltcnAjWFZn3mXWNo
oEtVHfehxSs6JyHfNp1DIoqedG0h58MnjsdeyU8cXb+YuVmUwVKPIOKkBYQ0IlyMjx9L9HalsdBI
h24pBdqVK6bWGNI5KGW7qI59pHeDhGyfH1pneiYcJRw5bdUxUt2grKX+6GgN0K62KYK7TK6UMETh
qm2fZbPMouwDOs48UcNl7Mav/Ru7CnwS7e63qv9oyldTupXd0L/QJunoivET4Q4g7dCnKDvsaO4O
FHqlIuQX/lm2/R3RJk06fC1aA2yhK3Jy2SI4IICF11FGDsAavfHNoyNpIENILPA001TQkWfkWmdo
/40UWze1AjLcZ6kY0qhmLEnOm2GSDyH8HwXVDb5rIs6BoQbf43onm5rpZoyMvCKIs1FfZeMFTbs2
O0fyCJ1HQVpfqKCyj9pSHmT5UNs70qd/oUSWIbKhxAGZvbJ4rZVnPAcRHG4HI9P9hy3oUuY3mZpz
P/fwpM/dzC0ufI29TJAb57mIkzx5y+nC+PEDOsdTEbDhVAW0VhM8A9eAdgqfoQ5moiOS5eHx7W41
nCujysXZ4Sk+fJVa4jzA4xCzDxbzhZsppGWhl8l9UJMvYSTaFyJNg8hwoAvCh2WkXWpTzzifFOEf
uVAHGYjiiKA5J/Yrfwd2YN8f0iy58NrUjd2ZKwkGxx5HeUcv8pNtbPDGHa4F715d8Z/shH7MXZNh
SR4RpWblIGBToHzsONUkDvx514fnAznQTf6kfHswCJv6A/Jm5/fff8C3fU1fWbKrrd2x13jjseKd
5HSCzey+21J/ZZfwh9w4deaFfVBBnXU3O20kimUezFKN+YtbygV8P9ieZzKqenc5HaqiU5/mdBEQ
KYpCAEle0yhoWxsLngnhQLuLPGc5fHClk1XDkIGOte41uSLgSjRhAy8DD4pShdJO9QhVh7tvpmNA
6stQ5qdSAZaI0dlXaDjdglrHTUSTckuQ20l7Uwq1oV0oh3Igho2wqCrRvNVOizChhItaM6ep+4y2
XgvgfEJ2INnAgZuwqmAXsqNawV5I8+O8m9RLBA2i1mfICmafpikzNUmFjpbZi6BqHrkzJkdaIwOO
5NSdWvMKP5V624yZJhjPSTjn3rWNHbFlcUwGUYV0z6XzwLmBxTlXHEz9ub6J9k+4anDIPxFyk4lX
8cTgdXdFS0nESe+ePz+0+mM2YBR2jlsX8alx5sboTJI0CU+L0tdmFwyRf7Ww7RQ8x8SThb94crRS
HrVfYJiqgwEg6uHr4dIgneNJkU96QDGUnJKz7SJenCZRlnzDHCDIsH7JGAzpiDXC2HduN+kfYQja
HlObldH1jfxDUv1/baEKSeDb26r74aoLVLa2LiQYY6nY4HB90rtukykm38jk7tYdqBDdgw51CRmY
YSeaxDbYg5YPB81w558knXl6O7CcIRPWzeYQCVkdCqezKDB3TSXNi13+8TT0vLRGfj2/RANRbWBS
NVtpAT+5JZbFP2Agcbd0hfzeYEwzwrcbDeSGFGxl6c/c8ViS0JZeOKpM9gHVNMvz2wvRfOjup0FQ
4kZ35Ksx2PFs1d5kptqQLbB2tZx2y08xanQBlvGR+IRD3W9xYhVYZdIxqRbDT2aE6wC5fAgtseSE
2tl1AwqebQJ3yNq7AoSH7KcUCJHQq8mNUyRdoPmRaBQhVk9m26mKOh/c1R/HZ5/XYC0z8nptYCJ8
eCXtZqtSfcHKPuqlzxqk14eXYMHikG5oLc06o3jDMY7QNLMUuuncuhnGk5lXayHOMol8i2MMYPBD
0b3DbXLrTGeGKLiTNiBRdTbhbPNLiQHvmA7wOAYhJ464IvAGHvzP4/4/4g9MbY7GfTTdhOacHigj
RRPk6UHCZBL6RWBCl7vmz6zzmAiPCMboM+3zfleUefmCyR8xt++U6z9/vDidlEpEGOT+oNKlet2A
zbKywc6Dyx+oLbspSVo5L2iY5OTFcNHiyGZaTZxmbJr1VhKGewvmlpGs5uv8d2vesfa4OlBhQz+C
7rMtT7SOPvWgrHSTX47wjdfUucG18jqWpnXnBkuB8wIetHDzLK4j12Wns5Ra11nxrCj6Z3Ej/ySO
SLg7fiOK9weMFkbthmpaTfCX1T8UTQoE2HuZx94oOUtPGHA2hf7Y5tCGXmgQOXku78LwlJ+yIfLT
Opk/X/rQa73UiIiL4lhv8oIx9ZeYaDR8yqdMqq1LU6tbywJ2SIdhgaTmgURiN6GKH+Ep9dn6zUNb
TPv237bzEJvGCInPlJmNCcYTPMPcNELMTrs5lI1fAa+G5okKjh+TGgRQ9NbLBUAaH7xk+IfT/Hvy
CbrVXVFiTyYuC690Z/GVbKk6tz43BxXv79WAYXFHfRDfkiBCRn2AdhnGaZbP6bygIcOxCzZyQyPo
bb/iV9kwUt9WQjNsadGvZcwSDaEPBeA48OfaQJ9q5D6yqY8r6p3npO4tuMLb3mrjs2o/ffkGv+wj
dZeAJQCqSWdeoaGRR6dbD4oxy6VJirI9rwqPgIT3A7sUHOzkUzFx4atDxEorbY1tmeirxtYkBPBo
iENstiiZ7evIQn2W38Dj9ksVmrmQMVbxr4p04Yb2WtG9r+OYgweZaUk+kSi9TjJXSNUtjqD1ZEuR
TO/oHhxviMV57zA/7jbWt+BmSbTP7qrslbhPkXGYSPxCVuxJzgEPzvVOVxz6YKaTCzfan+X7Xts6
owLl8Pk4Bw8v53xY7bAzAAOkZnkSZutseA5Uptm5CZCv0wdeXHxxRzX1X+Mz4trQtnSUrqPnwCsV
zG++Hzyvcns9qVE0/bBXB5qt6Q5aZKtmCAapkbqxeb1PJO9RwxvF4J9iFgzg4mGTTpKl3Pgul9w2
hKJE/hmzs3ZkYFpwcGQ3jPj29Rdgs27dUXbuwEhLUL4TLk0nl8K9dYKbldmoygGT14UwoQOVWSTg
LE/qUQBg0ciyRmcvMjb5ozmL6MA3Sj37F8ckCpRMuF8zk9Y99i04b5Drq65kwGA3t8VNSvENmPM4
+pVpU6PMhrpc9qtHdJc6AolfJWMuiSO2syoPyCrvKkxIBENI+pbRXh22o1NytO17qbMe0qbRU4x/
+WbETfDGGPmtEXdq6oMjXY/YdN7JvMqMcmbVEDtIz+/foQNvR4vKhDZNt6CUEMsmQh7ql6NlnmN/
3UGi2eYtinKLk9dgJXGTm0DhBYbrQD5rN3gYWzSlY3FZ9DcgSkFYMNSwMQA7kUo83Xi3psyjIl1k
m1wV+VRxO4WStMt69L1B+gCAG247pNpdqxcBVAxltBo4KKdDAonQrILTbPLzKKrQ6sRGtMQcIZDZ
VuRvV5GwUEYhJvPMHByFw2Ul4D3S5QGJ2iVKJxvcOhOrIHFklT4M3yjTi+R9kTcG6SqIm8lDpxwe
JYWT6D9ulBHe5TFLRuu/sA3qIHjXSKw7XFdJzDdWO8FCn/+h6KvejXlVq6cB6nzIA8lM8Or7VB/2
EScyZLAZ85D/SfcuXaF6dX9+g/QEtQOJUhcNAqe/l1kA0S09PNMheZh9OzIX6FqNvB8u8c+SpDtb
IGeULWLnrupXmRrHw9Plfcd8OvxIoOIKGIen4GOTTathfCybL5RM0ECCEXmbmm/h3eAwC4Rx6eqa
0nUWbF04APtQX6HIF09VYmOYJ3CaAsGGrwRXxT/HfAwwCrls16+/12bqc7o52LbbnP4vLDemZBP7
2Atajp51i7Jj4Cfw++XOV2BsExXfTc5Y2sV25tKLJJaAyxx/iBpBY5YVWoLCq16OK7+wmVOQPTo3
+Ff7I7Wg0kv05imyxzdQNimjWClDTPCqNzjOWF0DFhsPklFdXGKCyzv/MZSoUYjeIB7JM6E/QVBl
rigA83h7N/rCZJZJevCj3+vFX4TXPXQb8UNgs0EMI3p0HeuhooroWisz+Q033Lz/bu9NLfSVCG/2
bCrQVtlgkxHSu5BP+lxjSKHW8fdn6DfYz1JrEeHEkhdjcuwZ2k6hcHq3venM2M/DT/YU4Njs3Alj
FWGSMnbpr9oxO5OmO7Kzu4/vkWoANEPJE8rIfOklN9TkX4J5EOkEz6VHk1KTOKgE0M6Ftw4kvO3+
Gg3ugva7m5Q5tm4tqiRPhWfOUKcYwCy22DVw3hnc+AywMMrmP/xj67ktVag1xOH+8o8vxyBMuoWZ
TQ0zn2haa6iMk5xg0fDXu2eHfWcIp4+FWNBZRkJj1eEw4kAE/6jsX+L/pCki2BHcSoPflndds8Ge
j4mtzqFW7Ux4ACq4WarspeB6ylOt9j7gJ3LuzkoozSwFrVrMBAIcr78LFmACqZp2+gJ7BldNiiG/
4TcfcjZqCrMhzgilyafNxsEbKj9KsGG8kuipW+SI/GFy+mPUcA84yy6ei5RIPWlMAD9C8cS089pM
+GvNfOFDs3Ihrs3inOH/djFDeVwlYqZSuFAcRcXKBfOT8CWbYJQRYmUFIKHYV3Ff0tAqgbleANml
tNSOUD9AtWRJputkrzomqY0G+VcIjxWTaJqbxV+KmD9EP9AncM8AmMUEGOxQmmmlxvDI/nibtJ6c
SHRzKuk1QYI+jnvXz062jqJI1JtMHvPmMRQC7OyqDeNGVdez+eW1cKNnPH0wAVwrr1XlvV49aYTZ
ft9F8oVoyhgcOJlw2STtGZMQeKnrpgOao4dhlJerAxc1HhV1Zm/yi6LGZa0ROlFGC2q5OazGRvet
sckeP/QthM6IbmSyVJccnN2G0RclUMGdF1E5+EK9zHkeutYadVGViDngxUzcWyyZak7o2ap5GvcK
6cOWIUKxPqBTHJN8YzIhFt9nfOKK/TN5m1qI1zSUszyVPiGrjyPYmjZaw7E+clphdfP8r/vcIsPx
DMdbL8mmy1PEVE43XEOQwcjy8o0mwUjKg6VCorZkECDtCxalSWQltNBMtmtaDffLkKudLy76YjVX
vCVGHDGylQDYDSSUqejTiUx1pIkknrJN/zokXMypwVYlFLuUQLiOBbj68s03tqzkkxBwZDpnCUu7
VYDGQuBAJA4pfE8gMgJt7x3z9aLkgjgzx0C6xw6PBBdRz/8QOjdFarBtdHDLGdNt3/4t4w9zNbmh
c4PV7bdtTvJctCEqxkgBFvylXXJGH1EeiD1XidJd0fgcDWHm5lEWburCbc/1nvtBCzhjE+icu+o4
Uk7bBmo+LFnpbBawhvxI99QmV7tg/OyKDy7KVnJmkRFBQiD8qrPmTRzpF3+/TIq3A5pU1fH8/lSQ
8ULlXhOn1Qjnh4iJHIeVXQPZpanAuFGckt+lFQpiWBN03BnZvXrElQSj5Uvio02xCWRiFdgXMnOb
QyqiSPYu1ypF99TueYv0yFdSlLaos1uPET2iNCKfw3nkX+raPdN/MwHOgcELlrUMCk16QKuajmt7
s+r589yvW37Fl+GCDosOKPSgPhWAxRgr1gnHsb/CM8/MbqN3CD0l2ujEX6MC6Xv3bsvA3RWHQgkn
V/bfQrJ7FHqQlFAnos59ebybE0M9LZwYZMM2PoHsoDXKpUZP4cC5cTwwb7lDA0q8+6uBl47wQ6om
w1ub27ACbnp1HRrbGttqkOntGbZKluxu38HKPS77lunjz1z65L5LDPH9oTyJv/TO1RLTakyeaCUY
vIcKrTHstCn1TXii+jhhb1YhCwJqWeJ71XvOTgslvCdMWHC+csQCuDV42kcnoQ8umQEDYwOQO8uT
iAQN8RiPFd5wpwepTG8DA3mgbmE7tSuYrOGofCkbcD5/fguyx8QWU9nOAZsZ+ns1MiPTMn06Lt/1
ZtPh6iarnYibQxEyBHwxOi+16qj1q8hcksmpu9tta+VmGloA+kv8biN6HULFXvu7IGhHs5ZwkL9t
II5fSInXChoq57xDDE3LaIP0qikeu6rp9wXPQN/Y5GZFwrN+tCVegqBMmAQE3jt1nZwAt0MAuwvy
y6+M7oD3fdktxauUD/1s8M8Xd+ueXZw06whDFqtOod2UkzLCd93JRz3VQEmQWLhjQROBHUq1vOFs
77XGYrItJRIDpF8drZHXrKzGPRaAm0xv/A2gnjczeJR9O1+E6ythZ6Zg1yhRPE1BTCh1gBPCTebQ
HcOUVvejbHfgG8QTiPpvIo5PZKNGi1EwG007HuHaB2XgRkxA7aLrA5n6Wwixr86kUpGT8msUIwx9
Cw5QsXQ+Dk8jFD5mTy2NyA8FZ0+/0WbqbL84gliov+5iHVgTARbKEMjxXklazdXBL4b4i5VbBTA5
gTW64oA7sxS63dRihaA6j+B3f7Y7W8meU1Zy/Hu+85SmwIOoz6Ivn2VZ5+qZedRAgJ3qjYqdilL5
a7zShKfCGnFucS1Mp/m62CUXwO3HbJlDjWwz7U6y4ShX/N7zjWO3vPcAybwntfGIG2YHzRcDDaSl
Z3Ck+yVb84nO5g/ZxlUQoUmW2X6Kn/+FFSysAk5AWcAiLYnUWkU89LqjRFeCsTJhxtLOvxncZbJM
Z6eegz42MwOBDuFBcgOH22APksgKXpc1tEcXi7BmXHau1L8ey3H+lCF33z89aa3Z0EgrH+jkq0Dd
6nBdJFjiK5fB8IxgW6KeYau4rehtxOE13oeBgmRdwVAnqiwcWECjZfIA0oj4TX5emDFEn/rDtiNz
FW6hDgUMm2syIyT1gza0x2IfobhbUu6gUAbq0iFX+ts2oxqmTanriXBMjBErolmB7QGo1ABoIlKs
otei38RUTwpu4yWODy27mitIPZZ3yFnGkkih6ADzxnZLPvS2M/V0VXQPGLNxiUKt4QbNyUSA88Je
z+3IMrFp0eZUj7t39+i9sEpieNwUoUeZixFOsvNviLax4BcT1XoNHCdVaY7cBmMitXOM0jCcTEqW
MEQfMXs5OKilNxMAmd7H4wiKsLM4F0/Xa181WNrvQxOzOIZR+EOEN2FXUmkNCf+qBkDxPHov2PnX
yClXKTYd9MDg/pHZSuxIdd8BPD9YKwJ62YHGCDSoNI1DqRQBHG/IPcAvh9Ie0KMmXXglZirCw1cu
x1DnL5ly0YwJ0M5X1hdiznct9ccSawYTJNm/lYE2vnF3l/F5ZGD8Gl1fzYHYQE148VumAH2UHDl9
H4H0VBXMFe4IJeoMCMvdIO+ysf4xs2xLTqHkBfdCiiGbJZMakdo774BGCLmZI3h5gktz/rTh9hNC
bQPtH71sKInbxWvVG2Vzq5KOj+b0KnA3WEdbgLrD2rZXgXf2YhoyYW2zMMDL03761zBCU3b+nqgA
2A0NmtFafqw9FN0VSZfmRyy4aX+TdQ3LH04PKfUm0ld7XVImm/ZYbw1fPbtEe1iwJBF2u+YKhNpE
WVNUmbiNwfOCgtD6vY4GhoRI3NSNtOvOQ9uGlAv6+/rrAKTUprechv/6ZNmFOW0T7uT07bPg+Uqq
tlkvkv6OsFs7slon8c/YSilhO1FQEEK53cqiWMH0JZXz1V7JK9Z0Fv3mlRe/HaXijIcL94bigkct
ov5istIyryGO0tudUG013YXw86eR1gav2w4OVmRnVQc6GMA8qZ4tn97qva2jU09m6oFFgpPUyGJO
L9cyo31aZYqKaSF9OY3z7IMZcOL088KaO9rHv799Fq95/VYajOmK3MtD7KiY/ImboF11EHQKme7U
Bk4rG4x/E/7sWZzt43KlgNzGloA5KvWYHsSBsg2VJaqmndv/6/8FPCLCG8FtWEmdDQ/YuvW0VUln
kH3DfMITldwcNHIlkrLbbCtKTsfVrCYPrret31BXo6Oi8SELYSG62X8QT+ZJ+0yRj7KxvK1qtf62
JC0W/Drqnxdpjv4NHgLWGwXGWWA5j8/lqWB9YBJbjYVFtkgKtSY9twcLaSzeI/gHS3SVJgTlbTSK
7/cvzuW7pSuEGxbxRmxyDRNDJiy/EJ+iNzex6k5cudCDZ2oN5wuzOF8WgRq9pPFzndayQcidrGAU
PsccBZQ4pmp+gceNdr0IPfV7g0hSHBG5I3py1ehvyuOjT5Fa3AivFhCFClOr4+5ccK1hkKnw/h1F
dtKNl5DJTs6JQ7dkbl8UMPZGfTRn6nykOdHhD81lE58j1B44Dd0wl+lSzBuKA41rv28wF5tQbQtu
UIFRXYq+W4SVnC3r7ZgVYP28D4/C6O6+qR0QqSje6YqTLofUzTZq6emypWwc5GL/3ge+Bb5k6P28
UdCdd+0x9vR94pM+hD2oXkFOLyj5Old25yDWS9pg7DV9xz33A9D8/tzBJ3w7GAGWc3+xVAXTy3J7
oGQPLYadXOibgWpyRL7mMePtKiXyZkexRMN6AgsiSa0PytRIhhTLkoKwoHsS/0UnWwNBlO3tJYSI
0kXDBnsuIWFsxi19tYO3S94ocyBQTGUAsN1kps6d1FOTeqpooj3l0kkESayIkUKe1qacVSPwfjY7
o+mgtl0MPXLKv7MOz3ltAo/keRPtmCURuvqFsvuo2bSkeCWnhzuZI2VHcL9QbracU2vN8MWqpN5i
HkhcJM6aUPNhj8hdNgDSyFXdp3ktnCzEyvi/7ZK4qHk8KFJFJST7LJKscW5H7eIN3fjMwzimtGZl
267fhQIaKYKro0g/dNfysVmqbLedQ0S8BG49py0Abg/S1CVLKtHnHHMQ/kGeL5MhUCZRn8V4X26l
SGLQ+yw9MzCycCFFJfAcvhktZrrki37OCA2o6r9Ko0pdQ8TAcch1xx7wGEfXt+AiLjVJ6lUytfyP
nILE792kebGZccqepFTpq8fy7EkTYw7hefI1E51rlU19uT2n77BionnNrYIQ2WfmiHDZd9WTZtuf
dxZCkchzD/7rBtpWTuAc34qovlsQW3EMlo4+xHzSF6iMfkPqHOCyI6kfP08UlDtXg6RmBMdg1Pf3
tcscjk3Hb+Qq0hzidJGj67xaCBYLuS/D1ZxUC19ZScDK/LMl8xdXrFlUa08njyS8R8tVzQpcKDkV
VS3xTCkyhSUbjuf3ek6eOkLvl+Z2WOJbqyYurZG2pwZP/xGpN/BKmu4vjwhH0TthszJqe7fzbxMN
e3ZeALtqH5oRDgTfMebx1U1WTaLaJFGjFODyWFUPaZLegX/JWrjwkcqxldM8DJNIlbl6d3K/ZJ4U
6wJdkEpJMZNpBX+cgtoNfuxjE8vlg35c47KZUi+VJtxxBslhS44qfgeTAVqPIpvxAdSDCuLFFPD1
ORH6saLIu2YCLGjTKhpKarsI8PMRMqlb1TwDiUT2HkIHy28jjr2dEcYs9SRZH2+RKs3P7kk0g6kv
SDGpNc91cAnBbGiRstDT7EPZxxqPJhQnIGvCdbOw2Vra3GKwKApV8XDwH+xJ2FE80jTVCuVmSQNq
ITyohPsMsbKmd3Zec6PmnjjKpWDyUACRU0zWYO5d8ggKWveEk9euRaRouxbtdOvuDHp3+fwaG0tb
Sq8uOEqCr9zwKSj0F9qyxwAAJoDeLNSxWfDyMbua2VEW8dVRcCY2I6j3yw+/9DXMKbuJnJFW0NWO
c4ogJkLSglKQGVxbrP+UTOhwGlzUh9qw+JVHnjJh1dH1Q/6FaW2BFXt2mxvHXysQKdj0W0mT++ME
QbJnMuyWgOSShymNU+IK6WiDr4p0m1XaHN4NYia3XizkRh+J6AFdlFQ9Ge53Awh7idvmhU17ur31
uURuMLBVs9fZGwfNB2wbaHtOYOlN/l9fqrcVrHXw+Bj1/Pz5CMO3zhCJdLMcxNJwM+Rl64eFvA/J
ffHAQpeNbcY/7L0rTcK5bWx3w3r3WvXCCAiFW/Y4vv3O4fe+JmuGeem854aRUm5DrLfjgqfRkxMl
BigpFENKZkuZsVqBvSTvwIqh+6W2asUENGAssL4ChxXBUN0Yz2Cehcu7lEam7FM89RfirWx66ziv
4gjRHx9gSEw73valtKfcM+nL5tHXXnCOxzjWieZJbCk+UKntHBlLscuOPoaAjVQaqFA6F2mG7yIf
1jyDPXZ8zfXxsg2tyNpOb8la7roFYt5dgrt0Pp8pf4yHo2Ig6EM7JjR3nu1bATj48qHZA1oHR3fb
qCZy68v0PWzdBM5bGlAySQygqnetRwrOY6nCg6UU0Mcaa6cGBIR/dCVGR/o2uun7e0wNxOR3jgJL
SipUCAQBFz8wo3G96g1Q0ko9M9ynGoCRwHe8AE+36XQQl1O3JqdnZLDzhTnjJOPXsGvlPbWlH61o
t+MPaYkqiwWwn9sWvjrDaaY8MghEnhrzpqq4oK8euHaCc9H0RC4DuH9fN/cmxkQPz1PRXCn/slMC
LPMkpy9Wx9PaxAR72mivg+YiX/C1se7Me4bN8lwrs17KqhrghLKWTR//DAYTyLAMmVEWpOV+p4KR
yrR5JBxplTaiFzPIjdUejOfeaqej2acPndxayPsOnNCzRm/+FWpKMqW5zXD+F5CeeKksax0OOdhB
pHcpsroRZq9Hpguhuhxz1DznmSX2tjN+nlZyk3v9pZ66kugaJtL44MU84Nqkbt4kBxiNei4tUSG6
YOQJcv0OVMY8SqwN5Ohu9pJu65zJdlPll4lo947L/Eigz3V+uOBFAu3uZRrbU6kS/5wG3yeKgBO0
f5mc+AH7FyAT5wJ2plvx0h4NfHQwnf5xwICdmCQLYOy0tigB17At6YLBjfN6GKzOxq2keMcf+vkU
COOz9V31Q09jQVdepiQE3cy4y4NZL5Wzb2jKHdmeUWUNOT0C16OOmnuTO9RfivPj+TPdy+JZXWpx
w1XBSQEWuZ1rQwTdvOdN7PqdjHtrcmk8cPjTHn4MEE1fVIF8rJrhzoCyULCNzn1ie4eMZ6tkhJU7
u9i0dUIrUQyzkzPM+OnINSc3CGZ0UuxcSEKWZV2G9OLi+gybD8xsg+gDKEFz6KFgwTPtvOl1wu9g
p/t1b0Dpl7J/YUN0w97dwzha+iZJSMMginHDXcGjZiGvHH4Hco/t8m4ApIuyGaM2/bXB3dYLfJRq
t/vOD/nDF9wzllKofsjTRX0JBv86LcyNSukV+zhUrzo5MsHxhLu474uzmBUAQSeQgA6ZQltAhD1D
SxQbCkMsQ+e5C9+E14evJM4v115sQZYNXnDGx4A+GfpA7g6iWvpyV2PwyC+6LSKE8YeWZbX5/ltw
nsjyiX7sda2wK2+lPp12b6MOQxi5529NMGhIm/p1rStYNRtWoMcp0Md3xYkGFbt4odR0/b8GxHXz
hGSh/TjUxaOb6CuO8rbObhOSUvXUGdPeRlKfMZjdryFjyrsrtuhkqUl27sOFCz8cYrxEucRsgR7s
/pU1SXC7xXDAvUfPsOlOLlQmZr4TfY8pUazopaNAREFSLM1mMyWN9BRXjc9hFZ+SSWImur6CqrC7
lVicxysShBG18CVTLYFntm1CNXBOBIpETdQMFxImYn/kLrd0Tbmiu+xn93q7MrxHBIXhSkM3ZFtR
jo2C/49aj1bj2malz2BiVCkre+K85kvbOAy2ZBwMMtiOQcs1a9nSpByWnvIklsSbYJpGoPUFEEXP
8lfIA7dcA+iZ4p2BnrokGo85XxIpsBPV9n7FuDWPexmMNEDbnWDB0mTBoe2VtGD7CH4TA8JhD/tX
eWe9sctQsJvVKfCuqokB4vvhzayYydAaWQo4t7XrzsCkYQNHOj1qpODW/jk/uVPE0A8pC/HOuvHR
7jHBuTaeChkUSq4yVk+389Jbi5/cMlsl0JtzF4D308I9zRyxwYoPpaBFszaCLvCmKXu4Hc/FAVBd
rGaGjeod7m6Qelr96Gm6K8g5SRiw7SbhuRnREiNuONzNufIVsTFBu+ojao24dEPO8zsYeKNXi61T
C0R5ows6fM93gKdQg75PEwIbIncFR8GWWs8OvEXSxmUvizFkZRPSUt6vjwatCaZP4P014TG9zPBM
NoB2nXO5VLJnx19cqomQ3FtAu1GAcFuXTm2YdwwXF8WPXyDhTcI+VCrnOqQNfyg+VAc70NK/cCyQ
lGFkLyBlYGOEBm0wcUj0XblU4FvX+p5HfLphyCGcsIAsNAbA2psmt7X7pFjHdyxwfL7NINuJLjH7
4oluv8Cq/Hp+xtCzH2WgNTEdAJLdv7npLvAXLORa39Fc1Q0ve7MobRVnvh0pATAqLunXlhh+pwew
16c+OhibJjEAfGpHhYGu4YsaY1u0LtjsKTn4hN/U8FD7moRLD5n4NeqECyq2gzAGlka4bvrCdZDY
yaouR/j1kcucE2yrEVRG3PXa3MkJI3ZHIXPDDMSWPitLbDXzy1iq8l36EYxx66YoHpGuFnBCvR+X
s9BjTbsgBeLQvTguSpq+UQ4qQq7gvqfH3j8cRV+KFohLpT/lc403Z7UA2uJzlaJ3WdpDUK0yLzXL
DVOGmiKXAjI4ErFhY4FyCpgEJ75qxh/X2Y4ZUkDfOCfekAEfGrj1g63i0tsw1/WY0kCmkykEVnJG
WVnC5Y8KH2+z4Zcr70upL5kHD9elh/5IuRMnNCMeUYHhehKf9xtNrLPEKM6AbPJiGGqV50i9KWG3
If6Hn5qJpvPFFs55OumjB8gE7K9lhmydy1ZjWjLspxDU8pXE5qlGYycaMinQKseS7A52gOEsF3+Z
QU0qgCPjJTuyICvU+TuY4XhtVr2n5JfA5xjgoQdLIaRqQ7I/YdakaQH/cBB9ESpzD2vfg4qopntU
JZHofolgr653C5hUKaPcxaWkxPNra6bTLqqpOFakHq69TTPda0qSqDZ9dscg0XosN4SQRkHeEHVP
ZPIZB7QC/5oYnPl4+gcwjKo5Kclg8kNcJNDdthqGnsaUw8MEGeqXQloxF2/x44LCMln6uctBGLd5
CkglDTcym+KqIMXa0ZPidibkV/v9rcLBzm6y1nMG/hUW2FcCSPxPg1A0TMoKLrEdcL6sh4FjBpXy
fTMk+TafcBpUwSKdHpZWT/BGoINrFNKOkiU/jURxBzyZfPSr3chTrOVeAKpcoq6RuBlXrwYLbcWv
bhdfebWy2i2SWheE2h2ZHagmJsUR7+4eMIamJWA8zi9dp/BClZ9clNgLC3vRwI8cPv2JGe4PO88l
WmWPJ3y+dVpw2M1yhsxVaHJLfmKX95fQPKOdM2/MDynCrXXJatehCZGZXGyeeIbStNZgoakssz5H
1/x3a/4iclvtWDuig5GO1EYiEeJp+5yT8CLArnJ2Dnf0Q9f1SD1i4qLEPhxOEMOgG91GTDhaqxbg
yCQI/2vhjnxHcqf2Yd2Zw8I9L6GG7WU914GUy2st8K4aXzoSF+JsGrGoaGhYLIipYwb5ZAZTR7fU
RSCBkt4Y8/zYSsFZyyi1aZ+FDjXTocLvKYtJ3ZwhpkFNByQ3SWI9tavzLUtYZdQcSRVUjWgiKixN
mXJb3wiofhE55W5MOa7GEGeNZkZZzziLCUYFfxnz2c150JAvbUakwGcFG0xi2hAsCzuD9yc025G5
f2HiVMExwcRtCvh35RgPMR+Ke59mMGZyvEwi2owBCRRwZyNBsYol7ywH6S8qJa/+7C/tYRDpFafS
BLt+QC7+ejR3oGovKp/5GrYBVhHWROIFb3EoUQULVhhPVdKW+nCm7IYHfD15WnZLiQdi/qXps0li
yP0bRS5fM9zWOBOlvgItWG7RIb/YZtjSfjLiPn0XlPt5O1ownI4/F+SdNfnwHA3ttAGZg/yq03BU
55kNUL4FnJRPYOQwvNqg6v2wLpNnoL+m899ho8tf1/fOC2JDUY1YheMNvnOA2cvbmV7LhjlCDtAH
fTEsfTiV6MG9ZR375rhbg40hmilS0vyHFuieMlcHhzPec+impDtp+ELQ0PwnEhqkJ+MAGmWLtN/5
TIx+NL0/nFdV7IZcjXEHg6KtL/gHptuiWVYjByaIreRAiD1A/HzL9OCrZShrAXXPqQfkJ5KLeoxe
VMxW1M49LppbKaUjhlFaZ5KP6Nj+/+c4UqIqrnkoFlsto4uihV+5aY1duBRUmze+qPHYhwx+JKBq
zSuSOD1V5nMe4qMQb4/bn5HamPXcVATI7wFWNUw9akosY5oZlQEXU/Od5W5w4h6O9Q2xPECZqW8h
74ttuDdASwLSAn91CM4dF2zbYPZPUVCbpPSQ8TKr1NOlXTm/V8YSRs73ZdzyUFC4H5CLfy/kFvpQ
ku/JDhJ3gnQohcHrcNIgtcWl5CR+sanhZzwwmqviRIze8Aac8VtqcKuymnc4jPyOJ7EwHT1TrcPl
CeZhiKMPGIRqnT4r2W+uLtt9hz70j5jSxG2oIKcmEyX44NNvlYyakSKEI5Vo8Z97hpVmczAf/nw8
dTPL8I/2BvS1OyOYv0J9UDmVDmgpxsl9ai0gAKH55n2LnaRbqyiCsw3oNilsxk74uYhEAws7ni2e
H2E5qn6hCwCT8frtI73rjnN1rSJ4tF2zzDWgQhZRLjW6lSmWye/684h9phgYTGUFOVgdvrJaihbi
mc/kgGV/OCApZDCJ4ufMzoqHR0S0cWlJ1anHSqzM4+0rr+HWa28Fzty9uiH9TWRJFVYjnzkF9YLi
L7Lreo1kW9x20leWF4XvElzbCd39a7JIW5p+XBA4KU74qcEAjbZnhNNUiT4CsRrH648ZoJXQC8Tb
dpi4Wt9RX1RWJuSQOlimBSSmbBpn91WGRLBCbd8ATyro1rPLXdkGQj65w0KKRzR5Aoon63nlg4Zl
aysmlIApPz2oy34x5syt0EQ3h0u7nndWnTHeMVyNqSIrTf4G8U+5lx2lII7jVnFEsY0E846DjcEU
MqpFg4CjMt4wX5sgqmBJGIxVFHCRUgmFQpSpPUtvGjzKEDOfLBDSydFOrxAFdKPwxBf8az8SDVio
rSpcm2d7QeNLfM/x/rAqBR8KMuy2Oge9CEddvDg6/28o+JdsqIa1AjF9VeEwjPcMbzxu33frZttR
M35webCGuOTk4nl4ik8ssiSwcMHeLtALttUcKQuU4oaSoZnN48KKjQ3Gd7sc3yJCMxQ4wYiYrQFE
E9VijHu0LjLiRrC/wXJunmsCbO24GwGwkQqs4HgR1sJrQU527eAhGHUow7Vg2fOR4ky68s7T//yW
eLQc0SVAqz9gW+1YhZpeT1zLP+FVddLoa1BFXwi2gIR/LWfwnJtyTOXE+GKEOc0uTdpDkRRLSm7Q
DV/vS4hzqWisddA7bHcJAv5wuluFHBJh0CX+T2B4hUkP7tVI6Tu5fQ4JiKTb5t1+/GKW9eUaG7m6
DPGA8MxmLLndWcmPZlMGkeLUjUaBUgN5Ofr1Mu8GZDOqFTi3ortwWRD5VbK0NOoS46SJZmsx1DPb
tJ+4FOe/D9EYhxOgF5ehhTYKaTGOgy7waros7Zi/uSDiRniTgYK7Lwo5vyzjbaeE2eDoyZd7uHoN
yVmvuf8k0LQAPvHeimAQeaLy8tkuLVNpq/dslCNZwoRXsNPHn8uyrG4vRHzHvQUXfgTs1vq1miZi
tIC6zT208f7aHu72pybcNRxyTJanwNsSExbvyqDu86FPqcPWtyYbl0t99nhVF9a6NfuKlrsSnqXQ
loMEzkGpKNPa6g8QvqbvIfjaVXt9CmZ7CACssn1AqnwBilV/oZ3mVALRXYXPDzNRsfJQO59cmDnQ
QK5EYiap2wFbOHktLoOhfDPcIpceeVUNg3VZYJQBiu83XaLH4Jtym9daOJegOrKa2DIweCqKs19g
dInQC/nQg3+MIywmL7qkWX6r5JLAPuGGGy02CLksMYgmtLfrzg4fyBDY/HjAhoNQXSoyCDwG5tLv
KFf0wnkEFSyAtKO5uSfS5hOp2B0vuFW64BqXvq0Pg+NeLEuK7Z/RfpM7nYZgGDIgqNacnL4EikPI
oKg+ttAir/iULLIX7CYfUnIAuyzz6dIddnQ0JT1DUsWNaTcSoG+mMueCVW2cOZl6hQUXqDjUASmd
3vxAzV0N1CO049L/lUA8WZ+uIJWyPTwyq8EtsgPs3882kxoHdrB1ec4pXnO+PpGcGbZKc940z9Z/
BsrrAeBlGGlR8mN7cBLvOnfGTRnEilYqtYfYEhap0kIWfqKTtXXbTFFSJP81N9rYbTLqB355idOR
b/CpNNwJubIsWon1xKeSkR2zUK0KUrZ/X2GQJm2GtAVybVnDzryo/B5VZoFr+pJew2TIE/oENVjg
3x0CfIO7oodD7ILDWHfFAPGI6XrDLWeNTdE9dzcl+UYrqFMjTHllD8TFCNwy9ruSMAGUvXdCTRWq
L5ogbNnxdtLFn+mAiecsYAgi/p4BcyLIaf7giWaNYNe6LlL+zm9rlrq2nA4kKZmgBLL+Zfz0JUcV
1aGVDutB0lrtwe7jSVcGlgoqO8EqpD7Lmyj0TR9xmih5YxdNCS9uCftGLqWP3NLDynDniY30Xci+
xQ10YWJBZnSE1dsmZsCSsKYZjvqj0i8RVuXtb7hvHrBsDPVPT4e7Mo81FQiDAxhA1qXPxL+ABnpG
hUKi3twHhHw54mHTzOXq4DbWDWrNSobWsx8+jkWchdUh+JplCGTs4Vdh44snWQ3ZQODzH0jpFbON
8JtYdkRWkxbwIE9kEW0F82oseQ13SItA2MHJIR5nOKadPESUyBPGMZAgIbLjjxiVUumbTYl6oJW5
NaIGfs9bM1c3rVI9W6vpFcMm29FKMweD3gm1vQST1z2BI2/TCIDf8fwLA9js4hJCXAEAnMBZk0Q+
uRdtH4DLg9yT9kdeAaY9haEJ9cPwWzfB2VvN7gozU2WbWWNVCcWlph79NNJj+pM23ApVAjMzvJ1y
16Zu61epS1wvTcasAyBFIRO6qSDZAF/wGf8YcrzOk2xigvZML8tYIlzGHNtvsTb2+f1SNKgxrgXS
B6+gAY6uKec45NU3LkfwXqnMJQ30RHNeQ5w4XbZ3bA3vp4lgZoX2YxV45X3/Wml5v3wOvTLGIOry
1yzSWDibZNIqBaT0I+9TK/xiHJA02B5QCAKCZSm0BNGXtQlx23ff/wTzeSJ11U0EP60r0qlHMktD
YB/eSjdFLnbuCLWN0sj6N59Af9tjujiin8sS7cOPw/OfiX4oEkIesiH6ClM2MyFxA0KsQJtWS3kP
3shbg91QXems4hZAx7qDWfu5ZmX8jVi1beXhX6Gdw4lbqWf9kg1Jp8D9UOwfWROdx5YblDmK3W9B
go0zULAAr3TyIJl91mzUlc4m9DfGS5ZYHIwSd8WABK3/dTSSuTbuTvY9bBNgaW31DkPcQeEth7GJ
Kj/47wvp5ZG67R6u1ZkWWHUFiRv8Oo5tbE4vCMGwhYbar+6KMpPa6AuvnC746Q6MSqZkFaXZk9Yj
F69YFiUs0Em4ps9bc5uMrLa/G2RaejjlvX+6/lCN1DDeYS+RPmpl1wkVGUMdFk6C7+wwxhaWVca2
mVkUNhaPkrD0qhFhXzWfQQqu6RftlXPasLSDiAeAcuKUMv2zYLqQ3vLzEN/86uO465XkrsqXxJbM
MQjNPTUmJIFo5jYc8sOZSKPiOAUOM5g2HtNRh+IgDrKvjAdbyQ4GlrTbrZES9kRv/tecpijlI7h4
4UwdIBeXpVcLnr8qq4B8FoN1MN3tpMKCxZMsmeoCcCrDwhmwZ2C3A+HrFGvNaGNTlZM+clo+ZpVx
GISxcUDH0ESwYupuGui1RLq5yhqD2XLBHYmhHiuqI22QJVX7zpkdSDz6xGQPt/L2fzwzieGslfvL
wTFMmzdLECDwnmfpGvxAAmzxpf01IXczeUDtAZLtbcbfYZ+3gwCZscyzfZTsoK88vedwOxFggK01
ZlWX56+dxuQ/cltHl3qglw6eoqsLex3CyhVgyNlOHaIPjlmdRsICFsGb73jsgqbGcPFNAHsEodPc
HgB4WNKevanQJ9F7WFV5J6ylQELpk5i03XeWyywz4DgbgIMnuxK2qrLi7hqZnTXEuxdCuIsEpCWC
CgFlxd3T5uDPcH4ySn4lrM3nugLbrzgCtQ3SjP7Pi0DLrSbK51kIwL7de5BSP9LDp1vywmOOvA3K
NlMy9dfngsyQdHBozZPi6t0BDe0FhEiBmwLNQlgjawyQH76mgX9200bytGXo/lezxqq7cSHkxlub
Ka/dP+ukHpMA+TzTViCEWJpKqbDQHcdHNrYnePaFBWFK0K3s6kWVF9FsYcCpS/hdrwZ/ee1dW+LF
eNsA2YpQPQOVTGzxs398xJNtHenLoHN/kQ5zGOHfAhVJ/TDap5j9gcMQ4VC9tv0hAnOfQu+yJ4c3
Fuz8X3YCWwhaCZNrcfq6xw62n9m4vuFyTI1+JPXSCOKtuJ5Jn+BGxSZ5eAQG4NCwDZXtgqHFbsMV
oFrKPG4nH75fSZajHpGEn355DFm+jO8alylMHpmpPhifFNROTyBYB6fj9nkwSYX0jv/bfDMYLDnN
AQ2OP2fsEM4I884aX/BEQyUhC2QnQYmCbZ6Bv4LiCkC+w541FGp2ieac8NPPcO+rGKvNRUdbPXhV
BAclVtGYSNsgy0kZf6eVnfNVWz3MlyhtjxvMsD/tcleseBdGABLH6ZwQOzFMhtiChrXpz/6WKIdQ
TAdHTTfmmw1U1uuv43iLsZtk5ct53qbQQl6tVAfXu58IefHSDyGQ5atFshwXpIZ8b52y4grSMtEr
+6UhGzr77zALgmaagTxKUqtT7bm9bVHaO5JpANSXD6tbRJBotTYuEKuZqkllR/RzmabAkoTLsawz
AqpaeTSBKkpRALPzWDr6dN71lGwa4ldi3/HXy78Lbe0krqAwbGdfZSn8Btx6pEny96dCiDUL1lPD
I6VEgb7YToVY9Sz5sF3zKySCgjR9CWMXqpK+TNLXc7GZOP6wVw1FgCQ1QhUOMJ4/bn7qwI7MYMdt
GobqHD9vlAlX0krQnXNSItaCOypHXQVbec3X63pKXjnI6iqGtRbm0YJuOx7npdjWdSnFTvwXn718
2FBvHSpM6Kzw6EWBL0PutpUT0hKilGurOigDHrOPnMNQurabAkPhsZRakCmUOSt1zKE0cpn+8UDw
rb/BAX13VR9CWqBTfwCtKye45fTAxSXmINOcN8xSOyOOuNJ5rcZUGPSH8I9/p2Tq6+FD6u8HpWYI
14Vd3LuSeuyrEpDHMNCxWg+sxj1QxWWGWAw1T34HsZ92pctCXa3e+vSa8YFqk00ibp+DKO3KRtr2
+5YQnfDMUUzPhanhCB/MoueM/QQ25tmO1UhAmhQO4a+giI6SIJJYCLXV2U1ThixPHdD8hfKcMw/7
4Np7SI/ezcXJusoHVdeRJRoo8/Xez+jlgt+0utJ2aeUmqmrNlxNSTodVvrJCNsBauUm4sWCqPFrx
STyEyER0MA4H4L2lGUSNAHG9gf0OZ2XMdvp+g9a1TJHfjo4RGEOR39fX7o15xyZndbyprLZSfNxq
AhNsz6EAmMYXaDzueXbHcG3cU6NytFkqYV/OkSSjRfpDnwZOrJAKF+PwKXtIuvppfnHeZQWOjRD2
UHy+NZX9odzzP/vEE+zUSeRx83n4ezTfeyrZIVVEFbXW+GJ+38AW2kdHkEIM1U+hzdUfEP1aNm00
YwX4l7fDjg6zagJy0YWiKdEObV5rgyfeN9jXO7hZW7Sg1pIGKMcwQJOUiYuX9S5xefGIueDTxZbQ
739kZuiEVbKM1eFfRSLKhOgGpmZSDMUkUJIj0H5pJK3SourY5iQ2suQfDZlK/qmSkbTMvh4FFE8G
xN2MUZE7SptPr0LbWrKGU9P/1ioL0K9kD7RqUTmVPvmM8iUD4dZc/Z6+5rFmgha3QN/ccinWG08R
bZWTaXJhPc5NpGbrAMSMRduBR74FL3VWG3+bkNjUfUOVyy58m6y7H4pWkCrKSFvHk2I8FSvVDGEv
A6Nmm4qpRcsxadg2cnc8335SYFdTJjYdE1AMq7lDxVqhnPnGb4RygcXq0YVUXgZv7HtJ0bwYJSYx
RkAH9n+owidm+a59bA+roUrzV7ZboGswXsOpFlXr3Yf8MRaqXNX9GMzwP8Z3ZCwYHYBWLpkk3uLs
9pAnBcC2YiyYYXhsu4fWdNPOnoQGEE+wF69kDlxL1Dsol6Tx8zU8cADXnHATvW/1ifYRBh2zAkP+
VyZNzcU3lKyy87O9/J4+znyEPCSPQumej+sS7l1z0f+4+gT7leIficFl+MNwQGYV6KRPlRGKl57c
fZwG29N2sujZJ9PL5p9jMl4IvmLohI+EY6uHBF9gDik1xbSRvsvcr5yGfWGUNeU6XrpGNpqwdZAU
R3kK9+se/Hpl5gmD/11V997xrAGW8MCDaA9gXCSM5LMB/45iNxokXybShhxStScKkCC2RhTx0Ts2
V6MQyOnM5TvetkZF7y3UBsMqVUZwF8uG+Z1XrbPQV+3dQGwFfxuUP1k8bzIYvixAFhv+gDZHjeMW
sGa25JCzAGQDdoyrYdLunAKXgehOHlxi4m+kPutNF14aGqNhVXFrrVufvmb6WW/8bIZY7X9x/RZz
8xNoq47QzVcVj1FZm/jy1nukBwpZUsGUoLIFEJQu+YQOWLQeeyCP+QwLP5sqmcm2XSnLs5tdh9U7
uQiS3u5cHkXtS96r4mAfshJpVUGAevT3F9WuFCDriJFOtuu7cI9K4aiQP9R3cajMf9zqd/Rpe3hZ
xf1YL4yhtXdJGbRSSS4BXkhFm5HEctGIroRaRkp4c3inyYKVNWOk0DCEw0aGs+5eIvu6UbMjkkM4
dSjHXv/Cn8SKrc+11iwPSM90lKNECxHa/WHS64UOPDbmAUCUVpNRQnv+kNeu4eoQC1lWpYBdfGPb
YdZ6Xbjg3uR/Bi6yZblQchYPf+ikob0zWWOlh/DeJ2ZoctkKzO69vhyf7QOnBZ27RNrLVFgm1UNV
B3Kac4K6bISQNirtYlrW5KgPHYuL8iqroCT9bVMl6gbAhMkZkYk3ylj/FP+t4M7iLiqniUreEEDL
+oL3FXBPpphmUy00krsr2xzjWT+pt6dlCzzlt29XqyGjhLnHpn4HEleRvOgyc2l7JcL0Lg5S0mQj
oegj9eSefzBIwGUZTkC/qPi5u6fB1c4UfYNzk46SvfRQCheSA3dkomdOBLGCY0KxUBbHp3BKuXqM
C0FuX4pn7rKpd/kyjbfh/zrY0vTCtenYEyFVbWRZKBweRI4MwJxwi85zV98Nh9OnCirpJeAlxMsX
zQSfCCBM99rHxP/bBs7Z9a/pzhgSCU979L05sXQRdV9vSorgE9SXFU8SL18xOf56Q2r7BRUnS0Vb
yN/smWGS0JI/0kQvnBeSXvoUQ1NBztCAULQrIRX/q0JXMUnyY+ftnkOaAUGJCsDTDMXRoXHj5S12
eqlMLmXGDnPNku083FrMcX+SUg4Me10gdQ0p3sxioVZa7SPepnjRFIO8kzs5vWviWwG34ooukUPZ
kBKEkfa4M3enueKfx/Jh5jbCokwGAfZ8RjQXOdYcX59OrmBWA/EYIOMEz7YUUikGLRhK1EAGZjcO
iOVQnoRUaw+lGCzUlc2Mu72Pka0mAzj+5wa8x1101WCaHsyhvNBj4mmZWqiQ6PHbGP1RIrwKsjcG
pTly1liwbEG2lZAyMM+STsCPrHWKgfzm35SnqpXoIUXXKntWLQ2ncBxgnuj1GREBJetlcUyKnr0h
355gsahbzZrCw4Pkb9ZPHa5FL9DNWw+eOMG0UD9AtKQVeoE74Z6QHV0aekbzfzcVfLNgHabkwKac
MFFVGdGf8IrcHQAhcoMwPO3llBOMJglC4ZW8XCg7w7F5q5bkRRLT5p9JA1UBWi5kRT3VCmVZ+2Yj
CIpb06RkxVLt5hYRh6u8tdhVK6hXS5JGy8a3IEIUFEMO87klnihAO15tJLL3HVlCw3JismnuH39l
6i08xrBUwADY/NX3xVwP3x705KYCt+tPizSlppg95qSeS4FXyHw6ZPvgqMjxxYpwxmajOtGHwSIQ
nW2hvLLfLW7J3NDUJV4NIgLE+AqbvnSo6hDvjMVwKR3g2Vy22O0XzAckxVGkSoTG9C0WQB+anU9/
qaPhjpuL3FakUYc2h87zna6V4JqIhqwk3VEZc+neqlJ/4UK2BfCH74qdo0AVuL39+f91JTPd0Q4d
AvpKSxYkgr78A1ZM20fPfTzFeQoUbsicrepKGwGanPq/K3l6D3DtBIMpqCTj/Q5jxxzh4DV71S20
O7l23QaDNCTT6LemvmbFxAJSZClJai4ZL388DbQYmyGEx+H2ytht8hdSZMhpgcdUQ0Z2qfr2xijT
nV8v7G7zi2BDgOPVgop9z/Qm0E/fQMV5g0uJppDhJJyUocQV30Fa/pUrt5iyQc2KsHUE40gIOuaE
hVAYVRxw266Vb5u3AolHQNxRmAYMvY5YhUyK6JJJRka6cfUcXgWJeZZQkuvlADkbwgeBuYBex6ch
Uj/1iVBfCvlTbgUKIVlLvdHGeoZ78sI1p+X+/t+NA1WjwrUo3MrnosrzC17b3+ihfFgsvHYO+D2O
svN66/K9nS6SUmzizjnciDDAAFC8phZVkGv45H9bBjLvDiUNOg7WjLLn/T2fqpsOXUUFOUYD48Em
avDCpsWdFspwmo0Dz0zOIbnkd1i5LCiIfxLMDLJLVtuwccG6JhsOsxERwJ2Rs9p9kWznBRwqio+t
w/Wh/nG6J0mG17r5I1boh56x3biOFyfOTkqvIvLbpLdfpmSVno6VZVcMOcjYcKgsPFarzmDdG6xX
fIH9AF0Q6aPWDcKfX3FreuuqglglHp7a7tGJ+Q5oD5kU3gOD3IRgk9Mp43hqMj919whDrtAhO1t2
FCaMlo6WxrdXC/yp6xBpE62yomuCeCJlvq0BgNJiRgm1JvZfsRJy7VZZVhC4D5NA4zjCwJIvhHkL
x4lbqiYLJHZvkp2qgDN8kDMK+PEwgZ58hKS0AgT3W/nyI8YJ96U54WSMVaVW1IPm57VDiJ1Q+l7O
hisPVNhsobEfHFHMOB14RyHbChpshCa/5AOcX1sihZLlxwq73NVHYS/Wj9Vy8fKzT3sW/2ET0mLk
lLvFSgWIPeW14g0oUQpIQxtGRkQlxExuU0vlgLzKGIsP7twHj0aDbPWUKuzdsylaXHwn+jM4zGOX
8LkcL21+YZY0qL87iCDT0ItmWju5X7hfbPGSPaWhSetE3Cznm/Rz8UgngXUgDOwWFRjRkejHYgXq
aJzpFQyEoNXmeZaE20eI4AbrjiTkibVPE6k/i6rIHeprMYS6lfL/1Y16ccZPW7MrP/0UqznFBUOl
6Jpzh41ycxUWwE7pHuqIGieSGXfSwnEHJZUrM7HiYbfUDGYfbYvEcgvMqzrGLBjeqlIXp5K+TaOk
HYiNSYI+sMA519xJN1vBXXYbpHD/1UIcT/lkNsRFWGUatpdSyyLyDAnWGzX6VLlcuy2JlL8KpQwe
q1J1ef6rH7k0zBbVWX5Q91Jmm1KpHmw1/J166K8zbBWyveDzF2TQOa6hrI/FHL2ZgbEjD+nBzRSw
/zhEmjLaTLMFMUYKoGs8As5ZwZI5VN90he4W02I9K+502HDOC1j0ow9Y2qALyJA2UdmgXb/gTTH7
JvHx9+Ra0m6hagVtYPx4/ssD0vhX8XlwONcOvVBc/NgzyI+H22lLkPCHHgD04I9bCDWU4E2pzP1O
nFuSGc5bg3D+ycCKypPwHHNGqOtxygusN/DQILoxpiibnPY1BiUVd/2uJNvJ4cP+PsoVVHs81iy7
5kVWs79avYUmeB69vJFT7VgLNieHBGk5kw78LYzgEmEM//xrN/T8nSR4MHOjHQzC5sYXdCs/B/QJ
bgxWIB+em27hrGMnvngXuyqlW+tttgjzPPVFCKsnL7vNvhhDWOD1dRNoGLBnEULaw5RVh9KKPCwY
02qjszwJvH4RnoAVgyPnW3fq9LiFCR74a/wG9YBgQaGnWJ77L+Z6CGdf5EKx7ABY1uFDaADQTRzJ
hvLRbtBdRjEugXmKDNeCjvCr1NKOuytYPSSqIT7FDaWViwHbT4WV7z30Y2bZHd34b7IpLdfZxMv3
NCQEuSCabH/ddXeA22Cp4L6U9HLYh8ZEBLNYQ2ToSbwJAEQauA14U5WiZ0QZXqnFZvzwPmmBJRbY
AkVN/Wr/xfyF+/cFnL4cat96T7DaL4Y5RNd4OymsijiqyrxSLbpjlDo6XsHyY2xMtN8NRg1bqnIp
ylMzV4n7XHWPBvJOh2SsZb4WICVG7rXjFRTNfV+3xQW5VojLylV5hU3bmYR2IsL6/Zaj8KrlXspz
ceWTa+S2RVm6iuBC0Xj+aTwaNtP2nkV3RXBAWMV/f18kFf+ccKWqN/Y4Tk69jd7jpigCMRdTDFHq
wrTDKUZy+5zRbCWRP13hP+tUsboa5NuEzRW+ZqsmHBRLm1gLz5INntrWr4wc7nEicswJD+SkAB/b
yAXYwwG+P4ZQr2Aj1gjDvfdxC2VSqHzfhsJzUIFAb/H8GhjBBkbvZIse2CKJX6MnvrMTgswfBROz
AvvtViS8BldWQz3y3MGm7mi63tK4Tstrdk7v4ZXxsBAXn3pQLc4zSBNziHTrARbLCPqNNWkSjvcT
odOObKunKzLHJx5UrHDx4sPCzST8t+mFOlb/kOaAN2knHwFNgrEnck6eZdjBF5yt+Ramg6tEfngn
NAbKESCJo9aZXQ3b/8c1W6LNLrFrKtkghSQE5k79XjldMVuNW2ML8aiMVdKadUpNHu7sDNPzrNYq
xOySacmzUN8Ka9hiFZINC1DXEkHugUHw0uatQGj49zYnhBTqiFQUQv35WUBvwBFdNyiVXfJxUn5t
15btqnQFnNsn7Cmm7Bd954L3feZFZ3klPD6EsrI5KdJ6dw8CDmA1ccTr1jp18CE1phAi1uVRaFcX
TwnjlAtmaZIAu6noajUDi4Wzng5D74C2YUkL0AC/AJvNv1v4VTz2F7b8dhMNzQNI5XjVma4si4m+
wTemSADVlRh6/LSzxI/U4/aeCNDBz18MEbXsp403a/QcR7UZemg7vGeL0fZFulkClwG11Rb0R6/Z
RapdJsaWRZxYuRxEQv7Bblr/5KSwTR1tQaEuKGrZzji0ZNs5YkOzJ3+IymF7Qr/AC2Kqp0TN4dOn
5gUPLj9b9xK9pti7Z+roKM2wahAlrdNGsAhd4lh7I6wXUWS6Nk1zwDzBOroIGNgxL2/2oY1WtebE
xGpof1nNVuvIgwIiGi6gBmuyirQ2Y+qlSDMRbbCw2hb/F7CMKCJRIOT2QDFAZO7Zi1wpIVBxpkcV
QtLCtEpucKMYKFMiOkwAxL2f0YFytCrFJ7Y/WYTGifFEqTp9+EbbrBXMvXiuJGis2zXpv7gEibx3
/+HIheCiQxYZmo96i9sn3PTqeV0M2au3D1X0e6E5HvG77NJE44pcLOEKSv207c09zqLnS6+lg/Yn
7Kle8aXN+WLs2VyJdNRM/Y0k2RaFd4AyhfoerL0pVQoA3xbNQxsbYJpaZ8MvzUCK+z2qyAt31Aa2
UU40IRv1Kzv5tqbYjhTMLGjyZkAMWLreghO8JyaTU8/7V5GpzcIbaV0/My1s5SiKcqwjctIcwStP
6F/lmm8VzDxBeMiw9mRN6whMNIXyCqWTUTmYVPV90hyw+d9hez3UfZG1Yd+vPiHZls280oXTEpZq
NQRCizrsbNrOZV0iwM0sXsjGI4983+ONgWUb7/zUhgRNEeejWPKUy+pJCTelsCLLxvNFc49FPczC
RF5e6dnvhJWEw1ABmpNWvhQeRoq+7Prz20TbVFO3J/nx7LPtfYSTUn8cI5KuU5q+Dm3oU/1+zThx
jrYv7IevsdVjFFG3TPtJToqYFwWMtljHQQHchqE1pCPPdD0+k+f1XEtc+U8NFI21mMVwObZgzJAZ
WRhAtFwqTMogVztDZtp4+eVBs3btGtMlWSUbEmhHeXbSXqg07ezdgAq1canRygShcrr1r/YahFRY
gbz5IX8JKd11dpnSXZ/z6LM1l5TqrOp/ztKKrRKBwwA+/uaglvF0eJdHdrf6XvwtmVEd5kMaA5jj
yKZ2+MurZ1TAkhpVSeNFgoHIX9Wqa2vuKb5eT0Dd1NQbyvi9XbtBwOW7zc9t0/j0R2gVjLVP7Hmh
smEvwvukN5gcfeEA7VYv5XnX35LqYMHvhWDg/2qurcINwiUFkoIsrOKfMjTJt+lKr35OUTl9PJah
tK8hKmBFkybqGru4enNiMqcHoqNVyWZ3O9IZGdho4ilI8UFWs/isSx7z1OW1FVZBADiYkb6NZUIR
BzTbxSKHYRlClxlkpQJ1B2+fR0XPJpxfbYjdYB+8Dp7ymijVZ13h940Nuxb39s+Lfo81CaazAesl
JYgekT6a4vdeb/Tql124rkLvMCcanCwUXrJ9HG4xYe5cAa3MDb/caLkTzEHUfDmTsNaq1QWTBLp4
8A2mMepj+QynbC2REkL/npqTKfw+QaAP/qo2SuVNwMVWgd6n8636jl9+68vqgrz6bJ8y04Aj/K+y
m8nhdyuYdMYbwR12x3MvqbI/C1zo252KgPP4a/pBQ17W9EpQZjYaPST3h0pnQt9vPew9cp+bigQl
/FTuGc2BonFAEVl5J4V+nBbqSVo36i7b602MyMdFydhWDHKf5pH0XfEo0PAJFw2cElKfh99JFQMR
i6kNO+92ubKRQR2qMLe2ATCnOD2xHbisPUwm2qywahd+dSvvRiZFTyR1Y2QK1lQ8dKQWrOBvSED0
eFNcbJ3W/Aqk2t4Ach2nuo1Y+MjHYZXzoZp2WXMmXBfmRtZI6n9H574UdNSZn2X/mA0mObmiRbtN
sq0hV3aF6XODgRlAzHG9YyhIlDqu1dsTOqnKLlRNcLvMhpNOFNLL2q7Z3D3JpqYJOwLwVsUYMLxu
8YBQrWO6+Q0x2uy4PjBaQPq9HjRSU1TuYBas49b0uMlk3UYYiVmK7PJVzDkLigPxmiLnJATk3yoF
noyCaGLYIYkx6s7HJKrbozC81wVK0U8XQ2hEkddTqpdWfGVsR1zj73Z/Sdm3VlJppnvsy075OQ2e
brNGOrWyGNmog5Ap1X9Kwy+ayVTu4XVNGu7xMQQfiX0X7J8uOGrFnL9R8Btlx6QNvFDE0xbnyeOg
DYsk+hY+oZ4kc+rsoWWG+8xouMcdmMF/wnevXV4N8OVOuu9TpF80/OvATN6Q3vHoYAfyq1rmQWh+
sueB/rzc5ba69ZsPjCcM7OJc3WN5ba617PVWZf9FWPTIfsLAqQse8FnuiAw4DsoD6ElsqYTvLGM4
YyLhv9HbprgPwZzPDhCvAce3Fpj22U5dAPKajexN9Senqt73kRzcCM49w+0coAdB6zvw/AE9rKv3
HpXz3c/xVwABsOiUYgqthwwU9qvYd9aICUVREH0JaCYUp0KL0FdyMtoS3wNGatK+eas1Pbl44tX0
KkAf+v5tKuOM+4CA4XtFxspMf4waN39KmW73LUIReRDoZbtD1fIp0IA5fv0hLLX0pnBoWNMGeAnm
qFxclIVgk5uubiDaNtJitTsy2xRRptowIzu9VrBMuB8WM6makpdubZP5NuQDzlZp9Uk4wg7S5ibo
FzBwUw6z57X8mSrsC4tO82+3oHbvOQyr/abrjxq5drjJFRcTIDV0MJFIbqWIh9ioc42C7vpWJueQ
jkoKGFV/igOJ4JGFWp++QhwbgzP0iUfV+LDCfBSkT09KCIr/grTE1Gpzms2Xalt0SAS+V8SqRGFC
1w8io1dLadxFLrbG5JmZpo7cLOp21RYJSyyz4X7b5PX7fJoXXYWBQeNSImoVJQ/iYnTzy2gOcdjN
iH8r/rgPXSqBqv6tgtlh8PWFv/Qa5ktFqpbHL7gqD2XtHtPmVX81a712yXwxP483gphyj+Yn6JkW
LPDcFsWqYf4nJAvqVJsv9cJqrO48jDVBBIDQYPnc6rV5PdwWU5XmukbNiQIVMXA7b50uyG2zuCaG
VoqoR2hxsOhflkhbm4MdTbPST0t5GWbeK/2TRFXjGTsxGl4nuKsbIBdAlEIaZ2uuVOsj5QlSWOkH
20+1/L4cq06NLQwB9tg6gQiy9nga0Ui/uy01GSZK7oL5yPJB4xtykPvWo0obnNNb7Qw3KS6QHGuP
gxu4Z3sKsG86iy+sZ5JpcfWgD63eOTCNFBVb2ies5vncOC6VXob6tGyFVqi2SzwEZBCvOQX718lh
u6+hwp8VI1MBNWmGbq0AJd50cbLdFErrZyszQJcwJIZaof2DseCk3WqDkJxj7jawX4iXRaGtegFN
E2ncetuAbgeqceqbEPa9MPGrymOdeVkaEVD6KtNSyJaBhu2FeKvzB2+jLymRSyZZ6F2mwGoe+euO
AE2D0r5q/sPlmb2tRJYzj7BLjkPouuaVwxXz70Ro5GcX4uv4+4UpfADi5xwmGdd/aSdUsOyj78vH
S9hTVIb09oRdLH0rJQP2Y2yEECBpxivBGOnY4WsJKRk1TCSagq/Hr62YMVJRI2UFlgEKsiVozNAR
bmN7BsvJ2nrq0aA5kRjHKZGNPfEeORrxCauo+4nZYl1RGERNkcowQKXfK/SmTGXdvsu9YexOryo5
XivXQY7IZcgkJths9/22jlgAyVPllL0I0iJ8Lvbe5c4rmN6359TXdCHQ+fGoFQrhyk46ClRgElB/
KjFnqaQ0fKIh4GWImrXvlwj6ir85Y5lG367aJYy/Y0mpjVyxscwzbYCqJ88X3ltT6vgRUq2aieGZ
QgpvqRR/FhRYdSCb6qzpMJrJzdiYCeTBOhUVJ/BPoGcLwR2wSjb8MaByQ9IWCcSLZ6/OqRYWZUbf
OiseJVQxhVmdpTw7phc5yoVCnxmqi4xXCd3/iuAIt8p1gQK+kfQoE0ZnDmVwr5f8tzyQPPX/7XEV
Sy0pHXBsKoD/PrXryTtv9hG/aGh2Bgo4H4jIC2hNqKzOeeiZe2jrDinrbV22fPC6wQgut+jdgB7/
K/xKFDAUZ8HvO8Mkl7VnFPi3SchkoET72CR2mpzWRsU7SU9T42AnUW4W6r/KPVoeFjmTMa8Ow2qq
ZBsGDBWgJscXe66atKQKEj1S5PUxIRDK9vlJahG2i0N0frWxXtuGUU28BVmMUnXyODXp/SFvpQuh
EmxXKCalNNodr6GALXvtbGz8fUE/AM/BfKsHIE5yYOWuxjieJqGTuClXXw5l1ShqsJ5B/LolgvXS
Q9/SBLFmXrjbFPan1Fi2juvhabvDrXkxEvfuMctNP+81djYfyQ0GD5t+iLzQJ4an2lLZu9RjcIP6
zGRToi5T5+v6U4qrlt7rxCszCaZ6OBVo/6TAJy2krYuK9uwpJfK9ubPempmMeVd9MVvnMQPh1v4e
Vofg5wQx4MEnI1jU2b3HfO5KzDxjDUytTsDfMiKZndtNPvpeB22kcFMBgh2VFwM4pyJSgth3umlR
ceLzThJrEKAclIORxW39b0esIjDzAfHiAbbx5HD1xMAazUEhdJVntM7fuFqa1rQpAnh46uqfuSKl
j0W7QiOkA+VtfWp974QrtLrYrywM9sIK2a4s7nmLCyAaCDjaA1IN9X6WjPMx9LVXBTkaRUodkLJe
39OgKT+bj2LZN1pQPf5+tU26+xDXhaQ173X6TBs9mk/nfZcCrVwFEFoOBe8YmuGq2rmv3BBCfOMh
8wuMHgJBNKU81yPnisHFTnKeQ6e8wCMN/DQ/KeHwf4jmB/iWpNcAvA0gsrsC5zFw9X/7NoZIEqu7
sSkTHDVQTyLdn00pNSZjDD6ID3pK4GsksJ3HviNLF1tcJRhVLUFUSwTDKFaxzQt5jiZeM+jCPmmK
tKSBxmw2XFMEXjKZgdzEmRBuJb564c94boPzVFgg0Bb4eRDpLLshqu3Nd1jzCeY9UJ4+Ove25CAW
/M/qRSmXDwS6nRosgWW0aVUPXACkGwyqrcSbZnl9oAadbogqVOPo2TPx/sFmcPoLwjuNQPmqABey
XIqoTjKmtN7vA00rDxPH15CFqLhNXCe3DrNO5chqaPZYZ3lMb7GB5Xeq+P3SdaCv/h2GdbbOzH9Q
5cUDS5CWbnYEhp357ThLIZ9PIMBe2hpTrGPOJTj+JmcEj+eUXb5n1w5wZms2qXPnxVAI7nl9I/MD
w4h1Uf2GdRtLKk71ALjPzMxpguklouVo8vgN4HBaPOCvJ+UdWPwlGQ0Huir43pV7avRtQoAcneZm
PTf9Ph93I3oE3VRqjGGxQ897GLEYZFS/wrpTtleN95asq+VyL6zy3rJuF08C2ICr1E8hrdKpaLeF
VlUohRXDiE+OXNEY/M9/HzfE+aWYH3bvg5hOvuGTCRpdpxHJWOzbDNb4eZ3fNJS9q+4OR/2/c9LD
SB0Jpq41e00EXSc4SqMNg0N+re/8uhAUuPBxOIFS8kwBk8vNewXKvu8XWy4aHsU/J+T+2hd2Yjxc
GCfYVemZmHq944TVPCIRm7elomD1iXkLQbOvDL3CBnqb2sOeOw4wHMskI28vQ8tsAWiRC0OhkS5d
b2ifl53KTMACIoYDiwhwlqKNig2f7Raz3dSeJWARxSLtg7+9w/KZLnIH8cU0PVMLyrnjPWbL/3fY
rZ2B53zByG75gewg1EBSUiFCvj7C4VNyEuFP1/OOyqwGfRLt8bTwf1A1bESGdjdDQjeoxiqUd5FX
YQLu2weCEz8SdQC+eSWz+KwccFvNlcM2aevr/+T5PIaaqCq2Khr1YZbH05a3AyQx6kU2Me1+xc6f
NUh6BnPtiyKQTBx9b/ZFmMcizSom7QzDAhtAK9haI9AIFmo1JqxCRm/ADuWyklqj5qbmfJi7gopb
alqpT1mJrDtWIg7PkY65L/NOweJSA1NOfiw3R9R0SMTW+mDL52qO10OozR7uWoQ4hkRWlKuTbPzT
b/s9kamS15/rn4Iq7ovUJ+fd9X1d5bb5Q7L2HvkuckgPEHMU4Dio/LHtX2VqaHxmDc/OsBQ0ZMMx
RcV4P1amFVeF7tFTEd78OyedqzItfkKOiUMyaVhky3Bp8AxaagfLcendnfinOoarWD3fBS+k3MIW
P+zQyBQTA2eZZpMnEwu5KCpy6OO6Acf62+gktDo6PDq2ltfhnHdY6o9cpfbKYqKfIbgoYV/hoDZ6
P4QajS8tx/2OEbomiudo25eOJKNjzj2sb601gF9LoYyo6JcVduXjJg4FaaBbp0JieUQRtEJTNxyp
JqBnUwrK8lE1o/PGdAGcAV1ji0nJW03l/kjfStwWk6mCOOGrPp4i4ugkyn0xzgIpAvyOZrFbNBgx
PwiVgi0OawFR7AhLgVXntTs3VQn+wOpT3APPoQocBeprG/5YgMzAC6J8kwKt7f2dituoS61kVnLy
gjE1D87yN9hOE8SpDgkKA4a1iVWcqZaVxjs1tVs7ndHYC60ZXVCyXQHMJ2NPA1XmQZ5DiAVDJ1pR
hHiqE9vaxSZaX7SIEziGCZRHGGem82bEOedERd3sR+6vXeTkYFcyzysPL3nLR5Prt/y4iIT/+L/j
wc3W+cwgHQCu3Vn+uEItV3jvJ+OIrwuLMdzF7DvBGFxsbq281DdWF+aMYTYFSxCeh+PZT6xqrY0Z
hj1AI0gVkQ8gRJi45pc/+T/tvsKFsg4udKwvEzClfauSzWzg5yhDYIYnPfto2YdfqSFcnf5m99xb
6jqDhhZ+HSL5yAEJ7Dx4/m7GGBNcS6Ylut2LKQ5M1k+vyI2UtSbneHaXEOXXzveHx1jeerC1T5Km
aWHByNfpnWu5f/t+W8Dp/JUcTGlltoy0ZwQJv8RrV7nwaYMlAugQJfRJGp+Qvw7lRb7Ax9wdx8v3
jIhrimSGPrj/M3qBDGoKGiCllOj8rG5Gtr9yf7Uk/Pu+fxMn2PaKEzVa11mBKGgTRClVlWkwDV63
0Qvgdw4VH8M0MqwD7NCZmIL3oLfXWTLaGqLI9ZCsu7P1tucwRYNJWQiUEs32wMD9yjWtcXAQSZ2S
Gt+vrTfzVHtQwHGf9irr8aV6NkqCa6b2EaeV4mhpdWa6onj3RI0Q5sWmKnnSoQsebQYPmiVT3pu4
isuP4i4sXfG8oSpoEZGzt0JIJgJWIoC2WwMP7iX4tkHOkW86P70b9KMLeeLPOdBhtdDOUWdQmhrk
3NIbYxYbt908q0k38v7N7SvKXuna/1vmHi96tEwlkvf1UPERVgP/22RCp5fTIyaSkDOmNcy6DY3K
p53HLcw8qVJOqNvoBCdhYpaUnsUIwM4GWThTYwCQoe9nDvAgz0IV1HVZDf1mz8AWZwap1evHODxB
rFv1kAzYRtsiPk0Wt0FvWOrGQ+1JX6JdtQ6JZmtrZz94EX1zyNchoYefe24S3ft/mFoxUbCH+NDA
DOooOgq4S2WQE7TUXF5UB5vHQIZNDBgEAsvYNvnevafjbDQBz5GGlqysFipcyzDTJqHXXErCfX2P
1tS5yONJOY8jGyrQNC/3CG8dYrLdgfxNfk1BT6/jgLGjTZtCJstmuS8u2UAI9dRpMwvPT8wKxb+k
M3eOwe3lGONWyymBnFIdCBcWuY1a25FOMf/1HARA82oRPpDkmqW4jrUIMrGOUFbFG51zJUQhIy4+
wtnPmSwygBYKJepntvguC9ALlDjRKgXCoU5ji+rfOOWa8aiTrQrYtzaTUDCNg7bzSQ6AR/Y4+xEh
ibdSqBoBoTPdivtb4yxzQvl2U4jkeguDaGpHixcvC/Cld1LIQ87tZyvuAl7ms1dTpRhoBldFIQ4A
BHWNblMYUYneiLHc3baGig3tq09b1leXhpu963zED1w6b/ObAtsjgWkLGm1uneQNY/+1wC2uOrzT
AVlACXpNOJYsxcMfpAxqxM0WeOzFa/QhDDqiPFo8wMzJ3jJ9iWKpoiLswtblx07fxFBXIqvtTVPf
rB2ioxC4Xk5DnQ4YJ2Bqk4P9BHUvf6OWKojqRUEDEUNzoNhS3Hg69J5bOB7juKHm5mvjf07dyblA
NLo5FD22bapH23O4w2/Uu85RBattxZQUyx0a+QbpZ2o6MiFuKTBTY7pAhrNmA2r84S0Yn//c9zQd
ZanKaUyKNnVGXHmzWUkBYxaPsdE98I0edRF1E6fV4qhpufL72mYVz3P7t1+2lKljsC4lTXAgayjg
FZwTXUkK4W/rQ0CjeiEpZ5dliS/3pa86eS6v5jtsc1G+386NZYXHcXjGy2050+V4W+6rpKfdNQ+d
cYTmvG8ftdPyQ+3CgbaPb8BqQL1HeSJadCHXcZFcnsPhllUKm2Xm6WD+NxtF0Wp0/sLhKD86pVbV
OL1ILfK0KOSZIrezPnHwekqmpK0+zGrWr3LFkbRP8MQVUayo3+0XjKhvlq+K/YqbIl1GiWRgG0+Q
k9he1ZHPtCjxb2kUWqtEhU0DsyGQYys9wymJmH+oLTpwLqVE5a70hePCxUacXUR1GVeyaq/ZCzTI
E4nkrqLotE8zdZkg4vK8T4KI6ZJjeLQAl8ncAGoI2P0islgyeFPkqkxT8HmJx1/QsjBkITaFwXVP
gQJIQP/WlAPFZRzjJVtU+uATqn4VC0Ot9yBqjR1Vg3/08io0tD3kUWkr6gnjovT4n9c41fCZvI2J
AHB846IcPKPGMuqC3ecBMejGLkzMfxcZQcDedCHuoaRovlFqwNviaavMf/Qs0m3XCMUXvpwU/+Vk
i+1ymGQR/I2OyLphtHHlfocElWJqeWWlHnaks9bigIlc+EpgfC24rhd//5CqUxtocvnMlJHMCH8C
9AD1hA7s2zKSg7PMq1qRTPEDc1A2SH9tKP4/pCfp7n/bi15shZj2ueyyrTuYnylSpiYp7phOnCji
3AwuAWik5ZC7e1rEK969BDzGJj/WU4jb39fsC1YEw5oOyJm80YVPJ68PmY4gryA6FoHC3JeqspXP
7E7K6y066tM6TKPlYHd2rRBlUfjoZK4fc8ssBy6qiR8wqDPoOvdYTDXUIHuKCn55Ewqm5zYBvvc+
jGSdRhkvDVtOF8ZmvTPs343tIfyvXMmhUHHbR/tLgWYmsDBMHhfg5CEEG5gIQ8lnKEGfGH4hrmiJ
D2SAbp8tZXkblCekjmwEeUs4Ouo5SwGmOGc8MOMUthL4A7EiZ21pNrE4gq3pSesuWXm3B8uY1pnr
Nzx8HzvNRYujsk8esb/WTYUUYMVEeQ4IeUZ1On0dEIw7ptCox5pd8cCINlV3/Y6Vbl6SsKUoaFbO
GLRwBbdL5JBI6mfIR5RmyZDF2HJPI4qAg+FwDV5zNFdGqWpTKnKgL9vZxn9n64pGfma4AvfY9FOA
kbcsK91EwVYq5kBAkTbcs9w+Q1l5wsOgSbBvpwSvfAzq2x8WRnbRnVBtw/6CsckAqvc5O8SDKSLD
78Zuinz20Ee0e/Vf6Fl5Eb5pBSZ7cyTkZ1uN5eGfyNFbTsA/SPRsUkiS3IALNhJ0XbCB0tTMhEfj
eiL/ZMr+5YSYukQFc83TGQzJUptomtMIw67T1UbaDaLJkLdFo0gRgOJWnxycb1ao+R6Xnpkl79EK
XkiiFy2omPR4Gdv5GIYMpdIkaeJJIZmHyzRt1tsI+BguGFKxQ214Ohwjyw8PGCr7upkxTyrx3Brs
kcam/aqi2Mrxhd54l5EWjOO6DJlP3RvBLElW48VfqU7TnXQn9wuTEhDNzipzKPkA3ZzKKB5w/DXJ
n8g3kVyUFscRxJxRYMNJgo2QFUXRcvNdjCpteLLJLpYa3eQo7FIgAzUAKBIeyINHB6/RweZcyZE+
ZUiIDlpzJqRU+qiX5ezxaBpo/iVxL42po6NiMYTUQw0Cct17SAP0AR+AIg7ltpAHpu8MbAe+KaoK
wI8/PRy3aboJlD6tWLQjInPQh7zX2VibBAt1jF07r9YW2nGCNO8UEV+LVYAXGva3sezi10NpUc5w
r3BU+OG/7s712U+WO3x3YeE8MkPbUkY+OhmwV0lp3bgREANsoHT406ykiK3qEaXS1k7ftWi7D9l4
Qqmln+FapcvyHAEx15EUkRRBgPXaz/APClxIsGdn8+gGNOI0LhXIWgXcjkgW1HO5SRaRpDRp7saM
wS1TZ4n/oRM7zORuKuk3g6mlCBGSIFTL6duO98JrrVYYTj00DMvPMFGnJMPgVOu1yrVxgcM4FjcG
U+CAfDDz/IdnhrdbHmXsOJNElfBHjpZBmmSFwQpAER4l1o39RG4VReoWIi0CkVD2j8qrx4/JOeKR
j7iJKDmqeM9mlSlcdMOBIgYW+KHPqwAnio5ic3zpRaW4pksuYQ3zvjMD3JrN6WQT+C1zxr7tIOs0
4G3VSjc8Oef7SO5SGmZA66WKBGXjm81cKuY1ZWBcUKPMfvAV+A027oizngoVnONATWu6F+b2Z2Xj
JR9HDyL6IBS2a0LiWFFK+OHBtLO8o0mwo36/tzTkxfzdiNRLclE4AWSIh1khSqUJ91yLvgdu9r/r
vJDwtg1UDe97dDSVPISnccZzHUaj5T4h8Nwq4OkE4J8KJrgA98zvXL1c6HODTxJ+6yhMdgZcOYMS
Ns4kHiUCez0rWOWm1KJ0Vk3fzFwbC7k0ZbBhLnQSeMwWwJJvlEmfItPbWyLeNu73ppodBTAArrow
HwRWEjVhLmkdMEKlRlr9j6INdTDIujoIgw6L30DmPaP2nHr9z6FRP7+HOciqTYRfF1VY3FkjZ+oI
762DFOXtBIqG/iTAfAoF7TuvsV2ROaLgmHz0LVf/A+6qVRi9PHDtm0JoFsLECfTAKqTHmCDErLam
tZ/GI/CseVmKOgb8+lk7EU8D4d9HXnc4FEUHnG8d8PLNJVeVdqZJ8UIuJu2kxVBfZvzSuhxYP9Tl
KzFQS/FpVYkpbiJ22bSf9EBk+5BitrarGOBe/NO7ZhJTd3ILSinoqrpsfD2E0jJC1/pPZw053ByD
qyZBPTJD6OnfCXxkxflUTh+5+hyZbMCgnqNYCvOThFybzkpfFtTIp+Btg3OQutCVsX4jK3oDufEx
JzsWOUA1xBEgr62IMjFekRGY8bCi2ldPR6kMHaEAvd2DxL/+Llx1xDBPQtIL22ZJwNkKps55RsWY
kIS6gZ8aYl8tI10hGC0YSA3l/qIkJ9OdD5bPyrgmCjoTrHqjyzBajYS+9Zxt+K72rdAEype64Igr
o3SQY5LF2xfANMHHQB5lu3RLDNKsHIPbNFyFfi/Fpp0SfuUK8+2iqGFxkqgAybO+I/AzGc7y+gGI
d438yB4aQn6o6xBNk8E4x6mE9cWPA1SpMBNYimrIF6Fz8fyI1Y+98Fy31idzxp+cTbl2eGjfdshq
ZvT/usbFYKxU7TVJEBAmo2RD0Yz59HinE9jAtSFF3Eh/uj+NipMCz6I/h1k1HLbScQDHkn0xJ9/z
NnoklgqwEWgCzwWi6+nsbiHIQUiqBP8JOtUGdowWjm7114hPTCoOrqdax8zvosRmdoVz2vi5JylP
C+c5CZQ0/BPAON4Wzxzp71fcMGTlkZqr7m5M+AbCOMmqm1+fuMdowYULa9CNGWSAZ1tSMIHaBvLr
zZU9qmVxkuLJjYTQyruqecXZj0O+1vgKF/JMWgvePXxM7wRpja4yN6jSn8Lo9SsFCp4paa9PloXm
7EV7HuSiKjwJbGLVFprH5P4O4MY0kt9o9nEW17vQN/xRpyQQ76ZUsLPd6s0xm0pYV5Mee2avAzPL
PeamgQT7EPqTN2H7GG9ougHRVzl7oAU+TQXgaBVTa4wGqCJ6gzmy09R5XIzECFbi4uaH0ZPJweQG
MFOGDRs10ajuIM/jg/WQlp6q62Kz1kcxq1JV/+AIq6cPJ3b79k/v+dhwECKFsT36Jh4tKhVaGM8l
BcKNLNCBSX4F8qzFzOZ+NaXx9/7fjdkt+oe+XbOLi99Fw1ADPaIxZ/KRyWatx2je1mxbDCF5bEZQ
yHVTY3Wl2012BtsXVvS0HeAvMwFHtmTtBXXtnuQcZXpgJZJ0IrLCe+st6jGmIZ7w21R0eXhwwCWI
YORZVjKyKVEEbUZqpLJ/ZPP0tff3y6xgRfJtRU5d2Ht8913p0sbpBYn+lL/lh8hKGO6qQ67iLgLf
rLMuhESxrxOtzDqoomjZbAWiyhXXz/dI9/+rIpFnrJJ+ko8zvD47tjlXw2x+a1eZzoUuLo4TUHbB
QbHfWTJjJnhJbyAOOIMawaYBiFXpOWqzXHUYaJkBbpqmL0lB67jV90yReRoC602HdNkis7VjaTSe
lpdtxHP1rrdVQTgbpZtProoz9GkU30Pq3Tlqj6aLtbtseHxJD3HGpNGoXKLoUCyzOZKTD0/3EEMm
O/vSk3GpunSFswhy/eM70YoUdHQCwZ4h7grkuNJNY1bMYuOyefecAtum5xVAPWVnCLCL/bO9NAMB
f1vYF/0SUDxk7TtrBg9Bb7Q1FwyWzQfOY2jggdyAuDYo3ZdSdPIfR+X38y7VHWNWrtmTknB+TXQM
SfVjWGvdxLoMQPjK6W8roE1UxPa+onupUDKrD2Xe+Ra5/c+/Az+bxYLEIDLzVhcR3YnVRw9BZJ5Y
6g6VDXqrcTWlJCqUx9XH7+Urzp2NzWz+Mtstz2zyEg4W2DUHiH8Br/S25aJGI3PRod5+TWbJcDOU
JJLPtaQE0XC14emLY2A+7suCdGLlY560HiMNXQ8vq+Em/Ctk4L8QzAoIM3NVCTQzoRW2WQvoHql2
/HS+bEPtzS9IsgIIIStl558pVO0JPiyqKAGTB8rh4qtrTLEpE3byaoEEwTHHda0Vrp39aCuYWXkK
Z/WLfwcCVINoaxcApYtxyWCGZZ/l3uMZE9yso0LDPLweX41p+6eSePOquXqNRV3U6wJQT5APCArZ
DSmSS4Uyv1XkKL1t/nGd+tAse/Z46tWLBUC/b8cShpWBC1OozzTe1AZ7LMb/SpbI4DLA9wPceIkZ
hC2I+rhMHV2zTq4uKaLmPwwUwDuhqtt+CHseUHEC3cwiHP9C3tAoUpTVlbLyHpIoZRT3HjGt7tYW
ah8IM4L611ZZ+V+d1mQXoZu4SRM+Mr/qUWYx6ZX4R9g3NRpb1a7MwndGA9PFE6Wyan0BYXFq5uy1
5Ryqs191skLTKK95tm8SD0dp/1QWQbAmirfwgt6aYeHmxxb7sgT01o4l9rOmBPX0seELyF1e/TKr
noVhJzVuoaOeJ3kPRLMCKl3KcpcwJGNT1vM8aqfbUwgsdUdZc4hJfF9XXHQ3Hx8h75DGqAb/M7nm
PSl6u62NKjPIl61qGLMf4rVFOH23JtDTsnW3JFdW3ZJGqvZphmrTMrJ82XbkRvM4T82JA/RHv6gW
/pReCxi/LmcaRjzghYIgbcv8fdPXPjCGrbtbRO1dYmNV25cn4kEysk8kz9SR7rLIFPyz9UXZ8Rqh
+0ErEq6H1PRhXeLFmTWy8BTakEY8iQRZq3uQaVGNdIX4eH79JCvuooS5YOLdrso8+lHApzQU6jff
iu3ScV8DlZ2UGRrWpR+VTJi5zNL+yvcH4jiKEgwVBfLE0Ob6MPNYVIJqUrBgLXv2hWTD1n0kC4qX
v9bBV/ySKPxk3+YrjePFxzBjlsvA2dapKXSddL3/o1dLzZuGL64396KEhAM6oWVeSU1AQkTw/TJG
9l7rD/WGH7T4+Q80ZDUFdSahBBE7qEZ3TSSJuK3KCn9FNd3H0JAW3Glk1DyekYTlHbUV/MNUFeX3
+CSnwH9ofaA2A2z79cEt8x98JPsN9u3Bsm8Liei1x/WP6qy4AGGqgu8juzQJADVswV6FD9IILCRh
OYCMa4IlrFTfU+uAFxh4Xc190qA8gZ7wp2G4gaSF2LjWF7kCpWugE5Tq6BLQQhznslwlaBmsKhxv
TVU3T89Na3G0GA+ceJms+h+MvYltGp3PLfnz/S4gyEavdGdHAB7QuO+q8oxBPEhNmhkXeU0Oevwd
/0K8iO60LRC3Qe6lznjDhAKimM5+Q2CLJ8PRuscJ5ZroPam4+U1OL+rjfSA9jxAx/F68uh7BBv51
cYtBO6jerC6hAMw8uGrOYPn+H+3mOq0awiIv0/dpY2SDlxmVzzgdHCy3/mm5O8ayJYqmm+7kwQ0f
H04zxs+hHTXN+GdMthVz9SdQ0FbqoRjrV0tdvA6OqXqv4n7wzTFcMYkJnI8xrqQpzFog9Naq3FqN
N/f4eLHwD4CKhhbqLNDlxHUsAiCjCDoT6Dyphg6RC50Gy/bTGRll6jTtP9iujwHhB3IhxI3OqNJv
KlCiadmyXg+t2irX2352j2nRNWVaiXA7fz3g5wsH7NogSsi8inCqkIVK3EDcFA1+4+q54cO9LIWr
ktMtFw+7cnbs/wqBSIdHA8jwC2seDZ7qDSA1AhYGpetsaq19C4xEpkJSXNTgYyn+gFVTmJp7Zc/v
ARXiOmrBEwe6t6K/pL8lkh7Y9im/CR86LGntEcnfMo6kYxNZiKDxB4+wHuaeCVGLP0l9EEpoNvFM
s4N75CKeXC4QlBB9H92UWebCoFPA0hTXo8zNi52t4vR0tl3m4/Jc5zvXsE1t6c++xGToxZxthi+j
HAR0AcaT+K3Q/ssWNvhJQ9+5+2lFn0y/73Y4Xd+qN8XUldg8nxE/PepCp/L92ZLq+9Y0TBOldd86
6/iOvhZ9/wMKAtK06NCvkhr8LTlqoCyyZ/Whml14XXT2dgjkz8vUmVmBGJbbjfZGAMm343pRiQKi
3mXa/FBQ9glltmAWzNr1eJPIvgWq8ivoZIuv387mKFnZ61WUL40cIegv2tlzwI+E35iAScf6SYJS
ransKSpveWra4jR1/XfLICVItJdQPtuHxJGyZS96QC2r3uIIGyOL1YLAG5j6pM9ftcNKMEsEWbjL
UP24dHLUTFoRHzRaT+U8Aj67hwI9zGqzZ+KGxZTkzGE5Cn6k0OpQZD9X+ORvCapPoLlaaANKRD/1
kmkqWaQdmEi1ZAnDMxdHTdV7+cv/lfdcCivs3mRz9vOqoAE9XmZoK+KLMzaOG7I67u8wceVMqr0c
JyHnvbikfCikrXQY5o4P6Tgqc9BVLSEw7J6ZDfc/CoNGZMfEU9G/DtS5wzkli6i/TyT+H/6uPq+g
JiNVKWlFpZfZBal7SeqUFkq/qd4PYNpx/ZfFvStZ3EmAbpT/DYCL9YH7wa8k79aT0o9E5HvlLk86
+Z4kPWYugro0Z7v5LiSpijESJ6/tieHaD/dnnsjsLFds+rEfnZC2HFvjUO/IFUdNJWajTs/2TtXm
LT39jDa/KhLnWlIt9ieWjalil6IHO3oyXaasS5irxOhACJOWbe9R7tqS4QFFOPIoqEmBtZRYDtQD
aTr+Kv8OiEbrsubZujQE3LEIcNw6aFlZ2+cLdoHHkmRv6RleF8FWJ08RMji4xshLZj1mb7I3Imn5
xoV8wmMbQ0/q5iTZVP4Pi3NVyms2aiPypN3zWR5cE77l/WQRukxjdCqOgMe2T0cPc6Dh8lidIcKe
Fi3LxrbhiDYzbkvf/Ap0hpjxKX/wy4MAoJSfhDouLHuuIZY5OYHVGufP5iaYsSoBn8LKg6XrLwHd
E6Q7uUfl+ihTOXFcClaiEuOCf6hgTA9G4+aQNKf6h2gCQMQ1h8ErH4uyoR+28y2CQ0n0RbtXnqvB
Ih7D878FIOucjsQOoha3P4mGxEMTCyakRmcbtQyExye2Nujsynt1w2BZngAM2ARnxxj60yUxmxen
ccNsYCcm6w2QRCotR+Gb8fcx9i0rot5ao0RQGzcu00y1B3TefDo6ftBSk5UsRp1QID+xte94ncAy
bkdnY5UAdTzOdnLFZPLjAzMuYNZH/oa6RCuULloZQeBOeoJ1OeNeuvbKeRGup/dlUrfj6gdQ+ysy
L7dFGEX7UuyylOiyOM6G6D6ALdIOIGB989tQsoMgNgucckMexG5N6Gm0g715volKqVoDlXSjHDOF
E1LqndN6TOz5HXKnIpVOUkY3nhqgE0SXF6K7XRZ1RwINarvwly7BtEel2NiZ2HRb42D0r+HWsw86
MGP0frMj/4shMjbsjyJ2JQd4NJ9c1TW8rX+jXcjWwGwHcbf7aqoVQgOxEEW3qUNaxn0+4TCVWcYr
fwVlklxWOTgNrlgBWtWATLZKTTzUJBavc5OES4xp8dK46Si6ak9M1byRb2Pm6Ga+lylFCUDI0Sns
6D1Oe38Gcuj2SEZX3kie5V7hycNIaFS3PUexgb2uIyI1aiBUuSdGdfeZtZzllTwbWlCT/SAyqVGV
D1OsoE6oGViWx/JIzeW2z2VqpdDAkRA/VRqA3c1ftXKhYYp51yq7i0oaXTDzEYIfTaUNOrHLFrTj
WxQCl+cyNbYHK4Dn1T0XQI2HkrXjLna04tG+edpR8CF6bUEJyX2/io/+RmXOpFatu4kXb6OruZac
AON9GXV2trU4FrT/s/iaZexCTKVkr9aKJ6NIZgq/42vFp1J9Pgxi0iaUfeHtxR6OUJb5DqHTLLlb
7GPe6G765FhK5483NHgasFboEb7Wp8OXBaKwRp/k7xkwqDaPr5K3Khvz7Ii20Kq5ZgMyeYvbSbWz
I7qCPNR1JPddgCWZOVTig/9Zf6cro4omxhZV0GyqtZX5EuV8bLNJZOUSXTB5DXDdviRrIrOQCwGu
I29Zh3TqzOIJ7YCvRl23dm8K3RwSI9U+StY7FTfBavQRA5ba07Z7BR9C5Np0InYMVrr3VHm79bR0
On28k2Yf0eR28qWlMALDFJnOKnswX/kdYr8eC0bRNKZmw9NGIRAJ+JvlXisPhExrB3irI2WALlYU
H3rZv1P4IDsWqAel2kSadrQz6q3zI0yBUyqxTl4tzwxk3JDwbh8qvzOxYR5T7thzbyDTiQTwdPdk
t7F8mOUfTHV1bUm3+B1XFOslZ3k5STcUQZQSWe7m++QVBYPV4PXZKJIPy5MLz4PU+WHK4GoYwu4b
Vw60cDlO/O/QF/nPTXS/VgqeYViRPVP5et5+d4DQEcfUe/7tih+mNJlpmsVnD54PSQ+6m4eftope
qlyMnNTBCscBprRrjsnnMymETiJD+BX3Wk3Q8J2piRxf5VDaOiJTx0YhUVKovSTWTzIIsOVCIEiN
JXdy6qEvj3xydoND4AVHZzrbjlICSN6OcxO7X960vhNfWb8lIPPUZBbE/ej1SjgMllR2C54XxJja
4KvCA+YNJ6Rnm6CI6AbFLtwAf5MHE8fdRd6jI317TyE/BwhTN6znNKSe2A2itg1Lzq3ZtiO3Qnu9
SDTChTi9w3s7hAUhLbUSZ2OLpVSb9oH0b6Sy5SOLyQdFe/5Ii9FwAmeKXGCOuMrJbCffsRRczxmw
Bt4lt/axDdKyEv1lCbIY7lj7vPjrGY1FZyfAOMtbzvasGfYKWa0Kv6efvFEVGmiAapK3ZX765JLc
lUiX4TZSizATM/UgZD/UNl3iC/7Z2GW1AQpErGUuUAp48V+bnjJ6avtLVz6YzUAV5eX422RH9A6g
IdvfYE8NChlGH0UM/dH4P7BQlvKwsbGcfM3dmAceZI3Cty8CzWV1r+zKrwDPyA3U0jj6qe69Rw5p
i+QPz9XHTgMSfXNguKivRQwu9faXSS3OGlut70POo9Dzy5CELqubFDi5dWqNFg1GDUqB2RJ3nSKK
O+eTIfIvShknFvm9EFodOiLmmIWoVCrGZRVjP5RAi5DfQGgHxyKbzb01lNmiDuPhRSitxV0AzmOb
WqmKXxML5/XxbXJwhgu216BTNAIbH4IalcLdPIsmZki0Zi+rdEMA5QEF9nHryQ9ZnqFriEmn2uam
R3dXS1I+kgBlR4NiCILnqgEQwtRWqpy5PF4TnWLmYlAHFLMdJEq4944SUKF3nVzocf7ib0ssd08W
ZUMncn89Ld1mcCiOLFZgvniPOQ3EV2vVqhcT1JO56MMZP4eUgJ2pzNmvLfetdNwBVBsGxMm/gwRp
X18HpfWGaVbMLzpqNuK9kFdUguk1QcCi3iqvZ6MHJxze87S9nsx/ElQ6x6vIITdq31DHrz6X+5Bf
KS3fR9FfTEFeB+IVzm7AEdRSoOe5XE49zykb0Z7yj9Y0ElGZaXvfpJ3qrpD6zwUMGUH1TRKEVvhR
IHW7NdbfflqzH9wtFY76OrwvMxvnD2rIie0ogtesPhuf8R4f8usVgky9Je+po2XgF/E6oDNqyVEh
7Qnr5bhZaAU4RFSe4iW58QLJ8HkCsyDAvVYm7tN0FixBFUV+NSwFgNLh3u5MgBwpyZM4pn/FTkkf
l4778EJVN7AYSo41CsYKACztbZ5IfE+DlLyfcSD+22A5sjeay8r7cryNjE0W66fJGorOFp1tCudK
HvTulpp7GOD1z32uPZpRLSt2gvDGsQw2DnI1rs68GYQbwm0T4+RLHcyId9hlEAyNAtHHiiVNaX0r
eKg4VnkKi+YRQp7J3m3Et4ZYkelzilaLGzxzBEhgbLww5ExnMh9+KXcewI3hLWLwqELoxNo4SZSZ
nuInNz47cb7Uw7cJ9sF57dFbRy0jzSnWjx1QL74Yd/v0MxjCaDMi9rW+mC9ZI2n5YEyIXAuL6Mqx
c38U0Qfsh4TzXuAbcb08L6uueuskVO5I8Ir2uGpCcmA9FpeXxGpXGyeJs8CTc32ZOTNWQ+e8z+5A
HziUQi7QxUSnVosBTGN+psj/OE94BPiNesWfdBFu8tKrejUq9ernZTdn6Jsm/p5hVCITNRx4Vo9z
hdTJUK5CtJ9ZJKMZUkQY+PSMj8bokBcHl65TWRe48V6P7ZV0T2WtbjJZbOq1t/BGX4rV6fm+5Imh
66AQ9RirkYtYg/OeJPOE7nBGc8btiWCiBOiYCr3GJAAhpU9dIgzZ6P6oL1rXVg40hR9uunQpddTA
OH63jyqUTKBji96CpB4bwvAl8FaqHH/7qsGHwtzQCMX0f9DS0+1HFp1v1n+h5xquoYIcFdi0dES5
AKMuVeLdUO8nCf91+LKVtiFVn2+UOAKUa00BTl/t61/tzRpWxlZ9gydcn2q5OGfOPQ3xXlBhPakT
+7FDj7bONTFhZItUk37S/7FT03V3CdBgykzUuWTtYpf6dGLKhmRYBHM7NonTVLbwFtgynfMjzeqF
5glUTBvkwkZlYPGf6/BeS9FsFgSF1nXg5rjH0VfSB7dxm37zDh09naD+J2jr/kJ0m8+3PzsOcWEV
wlXNs/NufHdDDPcfDhUHTFUvW61g9kh7kGOo+cZPBBkJxH1yzGV+43p18I1kaotuMFoh0EAFizYu
yLkEyfqhnwnakpKoCREEH+NSNcYIi5yLqoioGLqow+yJfuYQz64/Qe2hyIYF43N3io8xA/bH21d5
7SMXQ8UvYipNJ0Xz7XGfWRMhhXZ9ci+gQIvcuJ2JZ+AEaUeGXV4D0aPcOZP3qZ1BhFMPFPKC9ZG+
72t9Gw+bysQom0VLTFKFVvMUB/VhJvTq7CbiCeTY0ec1s7EvuoAti7fiXUjnYDAK6deOB+EGANF3
qxrscVNG+C3BZJ2/7vFYPuvZxNpT2HsFWt2Pt/gZzH279FSK0I8NDpBvQYf1u/bCO/rec2mgUI8Z
O+1R3wa82ePEvUzh214TmjHxZOZLkt19zRDmoDST7cZl2RQVF9z+2CchIPN1Cwe1kN43gybo1HZh
UiNTVwZd05nspDkxb9Q1RqZsf67B2UgUKNa1OyEjLailL/uNbj/C6pLBwsUuuHI3uQ1sh5KiJF/i
vcoazQxD7Ttu/uftBnc0oWFdAvNsw2Nz5yRqu+E9RWSz7REeTXXvn5SvlQrg0Bjes09iGDAYLDBL
oKsfTHULwv50Jfd10dFMl4i+a9AapcQgpCvBGmkyjFOcw8h9u+ZaYY8G6+xmJ9cRKCEsiU5CpWp1
/CrsULjVG00DrKpdYJ4dz5VtU4j9AorsCqH4GIbh0EelHOeG9Uh/vnpIoM3NEvJNRiUv4DgQe/2d
+KMl3Zna6jWwXqkHGUWWUnWhvm7ud6n/O5znX6EFcKL4qiNYZFFjskWYid/v/ulH6IRGZrNZ+bBM
X3agHUJio4WTf04DTFKVU/CnK238f2YNMb664Sr87bYxti+if1IW9AJDGbhwyH19PUC7RO7si1uj
2aLH41GZ1kQzgIQh5Wd8Vh+F3OWrUA+RUV41Eh96LXObzz3ik7wJadX6JHhpgkfq6K9oSAvvw9kV
J3Df9q6JwClgB0o9kZ7sOCTLamTHvA1kcXmi4ybAhuzQRYeYVbJQb+LrVpGN9CsSmwHdYetWyFIu
3taAiZ9fXZI5fxwJXZde5Ul5YH6ej1bLEhkCXDFRLF1TuGiwLhZSH/gM02c08nQMHh0fMCM5QK3J
EhQgpfVlfvwJTO7dceBMmm6yY+4CBr35XQxOrQu2vjAC9YZ5MGU9zV+RVCdHxdHqWRE6ga1q4Og6
Gz1M5im5Zqe7Q7IXgn/AY3U5fssR6DrKeOy5ZHVfWjXCH6bkpB5nkCvNyaQCcNAreeCRsha28gvD
YwLtqlE9SPOZe7S/CHU/82BgT+ZmAqfvMscCqSXatcw1fS4ArHpIONkMMbDuyC0JcCMV4LLa24Ut
WKnK0Cum0/FkUPS4mULe0n+63trtRMsTmn9djZMN3vFL1APb4SMoxDxKekmokE5qSegrZgvid4rT
TOd7xPtFmyjvhHTwjPN+Du15KUT8fJxrN0SHKY3q1WsDTxHimLDqTRaGXTtqbD0xVOr1DxlaCW9Y
Bthtj2CN1V08jsRSkZLDuxf3eAQOq6ENUf6yu/piGX10t72RUkIn9kOYia3ssBP28Foq6SfskVju
KVIj0v08nBY6ly6pw9mINrElIew2mq10nf8nopws9yv2iJRC4SioAVgEKr+d50psnKzxfAiRyRlG
Ym4jO9PPIRGK0cy6XHJLswCs2Y+RoPvpShHMMXB8cH4+Qsivu/alMvAW03L85bHgOdVwJXFL180p
Qd0Gl+s2Y71pN+k+TFX8eHCwKyT1TYxg/sfCnTFAWHT/yfrgn+Cgdt7xuXtzESszqfDMKbAHmp2s
UQoT8R3UIvV1jvracn+h/ooY0YAk75+QXegPQelBSQChtBRhkhtxqpwaZfznTILsbZOFhjTezgFo
s3u+Zb/F7WlFLCDH6vs8I2r4vaiuYvEMdCy6yQKoeKiMq7Jl+N9prsNRz29RG+NC5fUd1GLin0dV
K/w89DE7TUt4NlwB5sTsuClpXWz4urEm/eiELW1PJ7+5lUD95J9ZbgbfPEY9OuiD3qAohrPlPGVV
zDFoooYebaTDPYPeOiidj1z+BcKTxwdIaUP41D5xBW2HsF9IlXcHzhPmsS6Vj3McMommI52EbEnW
a/7fnzroSr6lXG8onHMViXFzto5+8KjmPxlfvrL52NqVxLe1+OZJsE4eHpLKP/3UMalYaZxS8c93
ASVZcg7SPaNqfMUZRyfbPYxDO2WwUuil+1HudHcENm6oOE+qPxKbrJ3HwYdYgaF+GAvAZ16d/kP5
f47n0twOzR7NYa7rnYhEWfSOaE5504IDTqJ0M9Mql9F8uI36o9IboZzbTpMXaUci/FXKovT8jD6J
Y/RAqBNvKo6zrW6YMyk+Mv7Y1zLeggzc2oDFj3PFe6chsvXrmi3uwfqM7WRLEkDi1pvLez7zRW/m
Xp0EtCqXAI/d57I2zlDcA6PXBYrONyV2UlWgMO77F7bingbhmARGbGLo7e+VaQjg/aL5fgX9TQb+
CyKiwPgywKGP4Qww/ITZGSTE/cXz8HhxPK2Xvxf6rpHXpYdZJCJ4wcsuTp62Y8usr+xNxlcCZrRN
NbEvd6iCQ4YVVraXwLSW7uOwXSYCzuP0anoCzz7rpDbHZATJWYZ6fvHuG5uUxGhoUkmG3+4fLLuR
Ah+nbcfnGv9J2JqEV5HeavT1nvcU/NEh/EIuqb9ygFv4v1sVokQVLqr6SzQYFqt7lWNzEN+ItS0Q
owxWtsSiqFcKDNtxEwBiavGcUVRe5TBLeShibcxvXCtjs6z1BsSVbbXH8/tzluaaMsbYlGc9slEx
ZWSzWLjHI6d1Ccw4zaZ0lt4YGXfQcYc/o52bhodVUhpJ9HptVAVN91J1YIoQZrmfr3YOO+3rXchq
VAKDvy1BA9P97xAnnokLU3WN0V+f1igVaNrlh5XaOJFg9ewIkV7LXrt5cAkNxSJEqKsG04maocXF
ePXjHQt6vLzJnZeyLRS1zoNhRLx2vEdi2+PnF15JA+FuNeh3t/HlI9//hw825a9Qt9eVVZ9Ca2Wr
PsCz1nTvqjJdFnIsAod/p2Hq2PzwMCztcC309aOA8I5njqYpUGpwct+uvCyLhpQZUKYuUW5wbtUh
UFjlE1YJhhuAbOwPIo4kNCF95y0vuZcPBRqOH5MFKpHS2pSdHehC/rj3muy1fJITCJvO/JGmswqP
9yiYgeurxdK8wvszuv0tVBK9MfKWpBrNH9owep86pZhOIh1JJlQqIBk7G+I9B3zuKZley5uMnOHk
mI53O3pGLRjHh55lqJvIKsPU2BXRYc2RMlXEYGpdFB1DIwUkA3Z9+8GPu743beAtsWvcrvFw9yHF
Xu1qRsCGDqyuZGK8RYTiCzcRdubH60KU5FMGiUNDag+hfsiKhF1gRxHxrZvRYqK8df4+LmqoQp8q
rXVQjrG/TBAKwf99mmLRH47pD4duzS/DojxM+1MSO/Z3qh5MXrjZoCqjGGQ8W2zth7tVhrMj5jno
dR3qKa3KIBYJWQC8c3Kycq2acufX2YGAwAkC3iZeikcQYyD0GxHdkPuJ717L6Osq3Q1KQG8qJ5jZ
17FRDRMenLEJpuPtYPQCuU6NZ5G8avOSDQIwu5Txe8klKAfom5ms8gM/aa0fQl2VvQ0oyGgaXPVx
Qwt1IFZjhitkJe40/VjcaFjaMu513w+eRSIC1LDH9QFzspi12DC7rat+wwG42krvXploatblMNtH
dX6i4iZfgN1/bSe+k6taweHH8YEy2OQnz51L87vyhv/x5d6HAx21gE45jlHH+Mf3HyNFFt6PwMs8
MK8QY9gdDeE4Es0VUqQ8qavlz+8WcR0gndS/U9YN/KjxkEA+V2smYh4oyOJOtLQmdsNUTauIUHWS
hXEMSCaQJA2NOf+tZ9gqE4o6SRjE89085YmLA4IbPGPOMzHU1HPn8W/Uvn33wuAQfZRqx9rkaFxJ
Nal4ir/vjegGb4Qi81L07tk7gR+xqxdpbXZ0Z0nhgpr8g95c0/s8vhR8yoWXWJ9ByYbSnVzptgWk
dhdN3W7DDQlPIYzUKJcxGJSwBoTGPxQatS1kAizfbd72nJjk2vtZE5p/XGdljb/IJmMNIRSSdLqw
hd0f0IsYOEFVLpyW7P0EEMpqUwVIuPfSYFY+qmdYSDVcV13l7H746c2YJbr9kv+6EOpKvsxXGDPw
Z13xWJuDixxWgfMxVrlh2aKjHP91Cw8cUrK3GALC9wAJNat0dLv2XZcrj9kHOIo6GD66zkU9NlZ9
LUglLU5CoFVKMHUYpzPqCjNrmURjmB4/3HzKNFfT++PS0MtMHyJbGYuNHuX9LHC742K4MPiVdq6G
ovRVq78jd/dqwVN0WPsH6+oTkHOrjejFcTSt3bwB0f6kB3eh4xvRdr9HNq9u0asmItRSU8ChKC9A
woZWOz7pYLTqoEOQTbuSfjPxtgbm2LAkPPTEi80Mo+o72EPSfLip5aCYde1DA7pc624FTT+SIL5Q
78Kp4i3SgxrZSaeA1UzV5PecTCRBzoRwbF/lhDZWyavj0O/iOcRSJTWlpH5yF1IK2A0olikac/6x
h2YJ4AUl93D+bfLezzYscyN3nzflCXKk0VdAGJUN9tl4Zjxc4lgA+n1paG5EgEIAGckEGLX/XxEo
bYzLtt6TVqtEoMfPui8CsTJPdoP8OO9hp1MeQeRPCOEI/3KCHBIudx6AcGd3tW5Mee3/Pqqywd4o
v67691SNPlQOgNdvNoM7GNpIeBmqFtlJodK6+ROPN+KhzCjmXeqc3hZCO/Bp+QIKbXJ8dvRs2pzG
QrIAhr9PeN0lQXY7v8qIe+eGlHQYqlFhsm/QlCMZe/lrs2KWzaSeaSxTO2Ub2tD/FpZT9EbTC51Y
WH8BQa0s7U2kpXxbROwo02O7uEZ/YMn7/S+Gx6MsPSzCZq4YImnz7mud6TAtJf2jcXptCrcSHz0X
Ajee7llXXnYMVK1gEmf4UvbvGlWisVRVnNqwnzah7D/0eTQDXyJxuGsx6mY9LV1i7i9SdvX4Edb3
inJyOzZ0P/AvJofgwlacHKUGd6MHr/ZiI+TxkeGMpsFrFbL+PCNbKzJrOJjTAKgU4f1PzvRI4gnn
EC1QIlflMAw77i9J2TBH273bWrJ98j3ssYfkDthgYlVxfMT2jjVTk7MHTW3SD4gnFRU0mfCrDsOp
VTrDOdwb3cwMlgq6I7B8rQZewrLP/g7oqY0D2kSlM8wp0t9jdCyL7mWnvyqKrnOGphINRTWcRlHB
uCavsP7H73x53PrlGd1m+nLBPt+0vW4Yag5JgAZ3ZHFHNUz3nKuGPpPaYJDYEFYWsNsadnUkLiyq
Fjp2Cz7uyGYmtXtV62J5GOhOfFMOQYOau9sQjJJcT40l8WDAFotzXFxKhiLqAA7Y8O0fNErYr0c8
9fFAQC4ZK1aBmsdgl1fsKqIFXglYWCUimGKdlJ5X8hlMIR4G9K3wLJo0RlNPV6BwMVLlGiaSkdtR
XEoxMhNxjp1/nLS29ELR5b2o8thQNU2j9qy78e3ncwZmnzSW3HV3M4lqPG0U5jUIKRVeBiwt39uf
sNZRFQIb0yddy6VbF4Z+HKd0hYyLudksJXn4Ux11v42M/yjrBwwWIEcKqPMbTGF/0+GshwOXQI3z
JGmtxBK0yeidoUYRKt8RH+JPFL/vOHLyciJ3ST5+9Gm4ATboyYr4Fc7C1sLWPEBboM2sPOQBIvmi
cr4jaNqhI/x1UuVbMuYYmbv2T9+JIMUOuLogn8xOkY4F2MMYbNJlBlhknwCER7SN5DGtK+rnWqup
jRrRzlx2g/P5DLBJLhMVZyWcHzKUcuDstASW+d5K7PLJls+ahw3gaKg9xMSl5By+hjemFsIz87qv
FO0Dw1ToYbNDeVNgYxp4fo12QIo26uDk+AWO38uAJPv3+2nOKdmSmfQ6uSomys5FN0GpPHGwDnQv
unHXe4DC1eKIe8cyxhqjX9a+35pNL3hw9JjQFx6DSnBKidT2kndG/wjFfAH8KMIaPsF0Fnri7Y40
ESUuPjmLfVac7SCj0iUT9gXvBSTzruxlxUVs/4f7Yep0VZR8dU7yUPlrhBt8I/42FYqyylihsfF4
0s/1jZOX0Zpk7yng/9nMGvhMq/OjsUmFz+V020E6i9cnuJIFlu6+YFfD95xmwnQYg8NiDnNDNumG
mIBU/f9d8mchAE531jCc9XWdbnIN4UBZJIiM644PvmgHMq8JpBu/MVLWWcsxAtQ62sDqF35YgUw4
bXwOSJynKe/WRYEe9L0cT9zKC+RaH1Vi9/LL2h/NkdISmrAnxcy2sBK5ttuZJ0PiDQzpswXi4YdC
ae3YQxGHgS/gBlfue3fbIWerDgTYtd0V45aAA1hddP/ZXYv6EVU/UsNOYzKz/WSPy7oU1Zj7fVZi
uIzo5Q7Rqhxak54AF94mGFVzl7lUQ6b3RscPUUcKOeL1VesPjeW2E6gOZInWQUATVVNRya7R/cBD
sKo3tmjQ1bPDhvAM9vbQNksIIyhshIfEBY5Uj6pT0cyNkVMesXTlCRFTxWeHkuXUefHGkcMZeXDV
YjTGzawUGLicuFAie111C6GaUXWHyoDADZUWIy+UEoSHxPINExFikVc/s44ush0k0tkjUtJJc7VS
tpAQu498Hj+vDgBXknTd2j0SDLms9T+hy8u/nPuBH1lF864dCezXnr6G+TbeZRmDG7NpJStRWm2V
Dlu6U9gmk8K2B+VGmir7tNp6AE0GnhRyd9qGdoM7KyiU36xpqlv8wqkmdoBHGHjGORI5TRfytN3n
XRScN6lVgvKrh7Ho216OP9DgwhLN34u86OQ1hIqB+s7ziNiG/REkWYfMiRgB88JpzwfssvhyNWxD
OP7fdFAleAZCArNJ8/6Vng8EebAnYt7VzhyA3b1ExMjaYcFyt6uFf89yEal0WBwvVibhL+03HfcM
GAv3rwbd4uWZgUk25z24TKsrrIykfLYlZ/jJV6LSU02yCBsvVe5b24sJUMI7JfMn/YOz5fp4o5Vs
CVd2MaAwoRlttg6+7vc/VD0DHAdI99B26qc8l1LrAzugenY7XSo2VWYN7cwqOrUGpkBnK+dwulm+
IsEWdOIKIyE4ATDwYrRwcaCMgSCyGACQDRjcfklA6ylMofQykKuA3IS6Gzc18ElycK3/AP77ORcJ
2Qw+XY9oLSpY4xh+Amm6QYrqptlyXJqYIF4bhT2xbDdDT12Ry113GJbHAhYoUwZ88CnTmDsdfibU
uA8DlC8yQMyt1DSsgW8JFlz7w+rcP5BL+bSGQEvZBqEyHypmpkGGl8aNDViSla761iuxDSda2eU/
cHnwzbEPobgjKVInHgxFr/Fb/3ZjLouIww4758xc/+RDdTZViZ3xYb/vjzCnZTl2mzynJWx0CUUs
ANQ7YNFGLayoezU57vTPHvV5eeWDcUg/EKyfaH7uz/s3Rp4/tTBYZUA95+P2ynVGH6SFgOZGHuPO
fDzZIeYFVW3BgK2RDdwfb6HZAyEX5jIv4ZLQfQeme/wXmSqXI6JVQaSvY1/AD291INCLqzZWLfIZ
Vv2UXNpBugmmHr/CSc/a2gcEiKxSrKEdEkRJhxaaAVNjVBarVRMFRMkF/RLf7Zf6/wNGxX2zj8uq
+NBBq24cDWm+fF/F0yY+/aL0ksM2lS7hkM/WmV81bKQHkG6uoM8JIoU6uQuH+siAwpaW8T0Fg3we
knCf8TEwA25d8IO/GFzEwTPGyFQg4x/r2XSODGhK1uCHpDB9VX8cRqXwfXIr+CbuLb4EZdEkEyJp
SLF/w8HP00wMEu+b4gvRphLYgl1UALJCFI6PNKvZaoh5/clMlLuVpanS+vgizvAhIqkGXB4lZqVa
llOVB/GoXSi/tzw3bRRz8z2RVm2CVchLB29iDbZOfWyTXNR4vGdWS2QMGqigLE0l4N3UiG/0gIg3
fDbia51tU24Cin7vXumnBTHDXHKUfqYUVSWPsADeNbLkDA4QLFjPhSuAQDCrB+QAGFPSLwWLhEZh
cJopVCKY1LJMBlGD1s4JT2CpcVYK3NQGd08xKg+CjpCt2aJBnejSCocl74C/+59ac/HndvpKdl7W
LZ49GywMKtJerGELY3e8PNGHBZyDzXE/2exUGovqITBWUz6/kJ6SpsfmJ3+VpJAEJZOB1fHHrN2L
TE2hOw0IC1Oyiw01UIQiunLQNWDjwxfGFWUtbLcepbkF9orTvsSMREkSVu0ECcd2Sh2C8TEOoJ9f
VLnbKKMTMOpiP5JD4P6Ijldx+dL3gJ5xj1UouGt3Lsb0Q7SwjdzJ5H4WYcCWnPNCO7gAn6Id1NP2
BxzRqQSxfEtVptrO6WJthbQwrxsR4kGxeC+O8BZdN6jQJqI4JfITjLayXHenkbkjTAbvbd7j5hf+
xId1PE+cjKmpvVFjK+95AZrmu5+BCmmqcBflbyFld+EFiR5NwtqU2hp9QG784+RHyUV+K8ifvO4w
Od61/QirGSXn6iqb72VJabwmmCOh4xdp2FZrcQC3ipabAcea3nEtDtxdCnenaMhG5Lc8hmaHXc/d
Spm+qY8wDPlMxUUevqZfCNiian5UyG0C60zV966r6aY/7haiIxkFj3siXsPG4iQ5i2AYOCBP0bWV
6XAoWtbeDMIlWdtiF9CX0bWm/IJzTamEjXafXulU/ARzqHR8PPWaqnSAk83AYIXWUsuoxhtFYI3K
1qDSF4zPnVPDRJLYf5MU3glqAz1JTGRhQmE5HaZQ4oEGTNbT57+DBPvI2DgIQ+BCzs/C1bb2Snvw
rleRYaqbsQG1HZ9FhEilnoySFKYAjBaDUuYhaAgRitmdQZgGbWptkj3PzCVSMTXY7yg59ruKb5tt
kCDHz06Moe803ry5Jmt8DutM2R8Em+o703APSIaRbdXdfDa9UaKs9pE0vpqAWjvLk5SmilRkqrxF
DortR6CYLsQauzfc6MBrMj7HF3dGLoBJq3UiTnNdRzfGC+lUXn9J7YQxMmucoeANVfCZIUHH3l8a
U3pG4uLscDUZjOWGsCOE4dQrnLnO1g1vKnqiYIWuxf7DKmPfDe0iWUCyHXNoJdwzA9UuFnNxNnzL
GHlSNuWm/1IhjWDW17WyZyBDauWnl5IxFP4mH66DxkwjC+TYDv5ucuA9c1w+Dv+8tdWn28W8j8Q/
GilUyN84OFxu3fZysi2f5GY/Trn/U++s1RBwHaGIVDGNSLTtY44vjNpbfxGm6mMPp2epkNxUeD0F
6LUmospvBVm8f7YO7zDSHiH7tP2pYVSD2jufodXVo2OknuSf2BN+UBFj9hikRJZgJKYg4zZyFGec
hUSPB9tUPyMZwyPGLhs1VBdk2bYaOvMFTefSqQf4eJZihuU+OOTsh/whzOhuUFoGJxx+L2WK/p4Q
zUon2aevezNFSUHVG5Xlt8NYWFYnm99p9unozLQU06ZLnYfG5ruhKb0a2q7tsxlo6yd37jXvqYpl
BOBKD21Qo+f4hPWXQtN6x3VCUf9FEdXyB//SxTp4ElRJ+8Fj9WjtVcU3IEurQlNTyMbL2wJZu8z8
DwkVrW2M3yx3LgU3f93CteSF0nKetldO7hnUsiJNPXvrDMKB5+KXmN8utJRxp1dL39LZMQIhuGWQ
mVh3rGD8KA6Ze0bgm/LcT8ZPm9n+41VKCc/Teh5jwCGJRV+Bub3cfArPMH+3jjE/mZ20/sRuHUEi
r9tXdE4DME9GWWtgUpm+BSuVvEQGBDZiYVEghlUp1Qq4wq8v0AUHoUnqUk3wJLSDH0BGEH0sbSpu
tUhPs/Ci2GCLDX9Z9+24KxDxuIuaLLGew06HK2/+FJcSPmsqqJ1ProZuVem2RhG/MMkziwLKQh7+
1LFe8R1vA7tQuK7pofAk1NsZpE9A2j2Tj3ASuoZcfp2GjrP3vpd0uuDcnure+rS6cDORDu8txwb3
YvhqEz/dlIVndlwS2QXkgT7Ecq2EAhwviSh9hqyTxnXBATclUyUDoH2lEF2X1rH47CduWjwSaS4I
55LNkusuVeTGePi0KBV+rejdseLAH7IzYDDorRuX1mpCBKjEgzG+t1h/WBoo99OetJMk4QDZ2xTT
DRqxGDBrqL7ak+uqtXER7GUuBRbDKrJDSy7vvODpurN22mNLjI777zv5ojDbUkcOOoF8SfpAGvKD
kJYzfELM/jM0vWfJIKIoJ3JjuqdM/2iItJgpjTJKg28pG6ERx2/Y00gPexG2hz1UdQT0j0A4A751
jsvGnrvsPAAUA0xNiR5O33SBDMUkXtakoX/xtt+A2/HmpyJOpDhzHafpA03PQBT7kCji2RwI3C/v
VLxocVw80/6j5rE8Sfd002SkuVHHRYyaKltGSLQFSHjhc8GY1H9YVpAAhBbLvm/ZZ/tjL238AHaw
Guj4IkxCfrZdGxmqVJnss17F47I2nQDUBBIKO219TNmjX3r0JD02w2Mi3m/BUCsFjkWSptuqLaeX
5fWtFYaANdb9Fc1Sdd0zsw/RjRDs9425EEtZx2C1s87zSNx/zqRr+aiQ60tmL+CW/ATtkWuG7S7S
K2gtBbINMJl/VTLp/SltdjB+jzS+191CNi2bVIb1xZOAlC7RuBSF1ZOK+azEpxl808dYAY1yLIFJ
1EiPWNewFDJ7RUmNF85IhMAQ6/1GDTw/PMv/sJ3KH2Y1BuGM4i+oOq7R8TjvitpQHPa3jAzDL7Pi
/h8yZunF9OYefR8i665V3ykB5dcYwafivBDBFkSFJhnZgZUhuJnNOtL0swUXCJEysw6PojYxqA8e
uDyjDaQ3TC5T4r4xdPjF0qHBk7eoV8g6lwve5sVE4lWGxJJ1khU2TQZ1s2sy8e9GBe8MmCzQvudy
j+OXHz+jXXD46JhVY98syBofo4NvgWltMg8qXLiq4Zz89/yaKgZBTcxcbvuWMSUHA+Xynx5FPeuL
oIpkqG1rPFy74xskT2+fksaXnIVe3QO8JWYqmk8i+N2zGNJqg+8cGNsuFyRrfpT033qooDr45l7q
RF69mTYLMOJFEWKDk4rhIUveMlzm0Achho4zFlQzi1Ore7ONCsrPnTldMw6ZURP+vpcegZ6CVInz
LN04E0AITDW3PshSHjrtyQpxsdeoCzQsuux2xfzTJxSOvmmHei8PnGgDghDp3e1wK8DCarO+hEBa
Yofy/VmDO0UPda5WYyBCmtivf/FWZP5ntavFH02Tyrf1VdzpKgxcS7PJ1ErREvL4PINjgQg/csjR
MgCCGIX4p0Xwz8YokBrLwwF22uWCyztlHRT2I1Kv1viLWeL/xndpvq39drBEWS76nSOLedEPrF/7
55VYLUU/NSl+BcVE2y/7P//j7C6MEzRVGc2otn2k08b/hy8Tz4f04xMTLpGVHjzc84KbzUndupEw
te+eGiYXVAuGozp2oH8EM2X8UaC4iJm3Y5nu8578nd+hot2gGYUXA6gZ6mSV1M6C6thcLLbmW0YC
GnjIVB5yBZwqacVHkeMnN3yOJENQ5UIe1R4ySzMrdxyKCJSQPkqfTovKYMgmu4o+6wz+FyOGYFVr
+MvdfMVK3OddstoY9dbQ1R0vFWmRXPCnNn4z77qRr60O1Yfd4JdLK2OITcQNQlkPJ+sR6LcsV9eu
aXpvzvkGM5etmIv/stJN/XOF1zEacU2zCZ/0qyscI9vZWpHGWdJKKFjZhq+lhtp1boJVjLTbk3gc
/zRn5AeyoFj6mMcgSmSNa0j6XmaHq6zpQa5o3kck9ogAZglVuGvGxPOrRH4QaGFr2ILdj0bK3mUk
GSctyVy2FddAQiw2iYzaQLVNncMDgKjC8lQXpbbtp/dGpkGbrn8SkbshF1LBFouO8zA4w+eT+FS/
aYuCcfe0hBlOqg2TjRbSb0ChQUurQ5IG8CYumrgi3hJK7sp11DuGaALYGisfl4BD8qDASowm/C6c
Q8KIXJXhpHcImjNanZEi/q+/blGoE/RWUJqF2OMlQvOtX/LoWbiZufQBqvgldBjQSnTpZewbW20s
xScejr9n/2z5CtRZpjxRAAm3mJ57d7XXGIZvcDBM/2SWJwxMD2EFNVACADHN0efP4Szz72fn6dhq
/6YrGFwqgDoDlnl9nlHPetRK6neVK4qJlFlFx9oazYPj4InnzPxUKqxZ/HxsinWR3+IhykcVUWpK
oQCnWaYcpwZBNwthpYnbc3ndFxheky/lFPHrt52a7QvE8V3tQaffcpvBPfawIKxjQ0FrT87mLYNR
4IEJb7RkNs/rdoQRBd3qY/vZ49dDX0neOEE6iYEKKNQB/L/mO/wG0hqQTEz9FeUGa3wvUcFXjTyz
ziHe1ao8y+J/YxnV6e2gYDbV+bVy/ohm2iq5saMiSLVJIRjIwDR0sliQmAKwrTFIp5J0JXzbpcRe
jqUhJu0ZaPwEhib0pqpSWTNfxywl79k3Oj61iepdJK6LJ36WEtwoTTBxciooFclfKfZeiD8fE1Ed
CN22qlqNT4q0xnMqPDF+1bo4otdtYFVTTUba0FKhxuudzfs85u9Gt2qIF2AuWPlYQKa9X0lpfPJL
lq77XH5nTR9/yXi5XtkXiJLrqymTeUAtRDlCUNv2TufWczmPq4++JOlCOw2tSbEN7RUmMzLrZkQG
UjvEIhHmdUJMBs+Sgfyen3vIRZNRC0Ity9Aj1BFNJuTSO9yituJNbWfkrAayoknPdaisdOiz//8I
WXjRhEgEArsGvjdRTaJdqpPYJH9jBmIla7Esm7t9GOhV36yTNmgBW38cApoMbHtGMaaN+dpG6Qv+
74YSi/d7OaY+16SF4MFMlemCCfeUmI12FRF5tzZlHsRbVNMyKWSvc+sEHqb5tPuRAjVZAozuejFq
Y64+KwDCp5HqkT10E9HOq1L240+GYqF6Hxyxqj25aqnU2Fic9QM2BNCvKphEmpKQjbv8uLgxXSX6
y+gUNf28J0iwt2HqMcRwfvGqqHTKi0wS2QVytadnKUoiFD/49QuIN9xtjiTh1YQHFP8esp1Y9RLs
LZTu+RNL/iqBuLqI69wRgBfwH2R9KVbb6dW//YzgueVEK5uS30gqRJIR+i6irL5aoE0iXD6pUZ6n
Vh4H02Ihxt1+Zg+0bcl3Gevm6RTD6ALokLr/kYBVEzXVPpbQi83UOEkgyO1mRXqNnODYg+Syd/kv
lDY8uGT9NWR/zb6Ay58zcAgpmEvMqOv6qUYZoXI4+rewJt+m61l9YAtEH4ZlU12dNc5RW8HJti6h
HhoZK2Ple3YNy7+jHNf93JNH3VYiMAwjVGYUpglT24kgAnw86rADu8l09tSofulVjpWVIyxci+4N
N4Rp0pTymQbkLw6Y91qhynIPRZGKqXyEsyOyiK6celgVHMMk7S8HFsDRJ+DJ0uqRFMwLVdOiqDv/
6T+lgBrEocS69thGWXRsCcXEIthpRhz3EZD3k469AOKMIuqg0hul8DpPyL+HP+mnbW1rTDz1a3nF
+IGKlUIKDTtUMCUXPQ8J+tc6dehGLtx8EoBJwBac3ZEKy3dzmusTc2QclLSZzqJinfV0OITQumag
88ym2fd71LOTGsU5O4T3cyZyCV2jiucUMXWnzv5LsEGlHaHEb77pLqIT1vaVZI1VvMzI7rVbVIfJ
6M3Npvz3xe09bqSATBRkPNUWPN16uIAlYKJ+6o846+TFrrqxpL2w/XvcNgrFFIyJP5KQO6VSlvM3
j+gEguMwkX7ldXG2lQoZ0XJagNIOzHMvW7R/PtX/TW3TZ/fVo5rmcH/qRnplor6l4HLjwKXnzlCS
XA75UBUcJblZq2aOk2wU0ZsRY7J+5fHqFIh7K9AQwStxFVVbXF1dzO8Inv2jOpNGCIl0HCZ1XMTT
nwgpm/4tlPmL/VkLfpDfzccMF8qeudir13tYkbWNu8ws4Jd1GqR91hFAhebfj/SpHqhXGlIIyGXk
djT8E6mZPiS8h3lqr/VSspJmbSA3cygJBwIeLm2XTmlW/+tYBTaQR5sPrz3lVCuiPxEHu7XWOleI
biJOAsq6bdwD+HpQGwKGMwoGmtVcApB8boUDBOyC3egRR6ssSNZkq6AAxnRTR7MFnznYhyNIRMZu
j5mp1EUL9xJdtS7BzIpAFUIT3+sH6F/aaiApzE5vA26uqtDRpTWJ2O+bNDioY2jUgIz33fOaE/ZO
pJlmtUBlHdmBKMMyZAg51hogQC4oDX1pAaB6MHZLjIXJyLdPsM7SrF7xnm+4ajt1F1g3xgGqbb5P
Vxw0zutEHuJ6IPig5Ef2ekQBvRZ4FnQw3G0EY2+61f9fsfFN5bnYr/oxa/UyFOD08APnmMq9LSfQ
5CwQ30Qc2cr8zdZ+QGO/xNfWzdVe7V+ASFHsNo4KzG1PLT/cSuJPrV93loFwln7Q09ZMxyVnkLO5
JDuMlhF3JOsSevsun0SG3Cman1PdsMTQa6pR/RUdb2nUgXh3QZ1jPlN7D70SEHvM44uM2ao0hdG9
PX12QVJmhQVxATmInaSBZtik01T6v2tUMlmlTLw4j0MxTB42Xuu5ds+De6kPkfKWODgijOzFNLFC
EB+7mFco1TWY08uevJHIFm5KhW6lUerDkSFtrm0jV44ZaMoO7mu1e+lbEElrjdhx2mEyMwx+7Th0
Kjnj5TTnYH3PTtN60kN+yvdRBEs5mXVXLzNMTvOQLhaHeZeSYZ9yql1BmDGDxH5xRGO4C9aZhage
QfGUc49Ka3WT3HwmUO2ZVicFXs0H0DfTpanEWk/B5X7aL7U29fWhd6I8JHTHJ25KDRU20uLXdfGk
JKyG07Ecp8Dfr/fPBHiRQcaDgC+ZqlDm/o2oiKulh1fTF5JcRSyqhqdcDJREcy90Ttg8+jQRxiIZ
bN23sIgBevOgY6eMVkc3jXL3QSwjKN5viOiE2O8njm2Y/uLURpJLrov74Z5v/88wrTv6Iw8n4OVD
9HOS9r+GPpzPE6Qvp8gzCzPQSnsWvSulFPs3fByznfUncoeCLoKNop9IyF7cI/yLTEC8vj8p1OU3
TWszH66UfRzH8OXnya5vAcIbqTk/HV9HXvRwh2gHcmgeEXgl8nIPsE6ij8iqS2pkl4zLxKzAAsOZ
zoFNwal91P3HB6SQRVmlWFjjEuWHGbi1RI0MDAvucey3tGgtXbNbbG2m6j06OA6or8NwSeRdwTpV
Q6RU7HMnbgFU9AqWelKparBFmuggnJdw92ga5190RLiyRIOAIMralYMCII4zeR5A45S2XmaKqnlo
xI1t++9WxEIDLkE/IQSKhqWobYuOXj+zejoJ5HZ7YkZbR9U7gQfqd6RWbOJOLbdNlmhDA4aw00b7
+AVgvyhBjfmPlpi8aMhxtHf6BsgprUazW2oxQavt44cnji9vAtjmKduwRoqy4CA3VGid+Gu6Ce6D
0ypV5bqghIvUbgp9PJOlPpNBVmrduGEYT5wI/RNPuslAeQySEJ2Wk4UQgSI1C+kBPEicu5emvnF1
CWMroJBcCVfyWgFPtavcCaEZ4W6tIPUx37ggeSSqzdbuZRVP9/Z2CgVnm4DVQRDESjv7lGdTICJW
d4rXi4pFi3b4Wg+AaMQUh9cNZmj2jwq5dMPFnNjcRp1G5ROj+pcjy6OdouT3YeejNm2PCbKSrNiT
2f1FdI+71C2+zMBErA6cD3tnAKFHVzHNr3pyFalkokZYinm3lnzYQJGek8wNNGbyGw+jRTFNN0Ld
YMNJ/r1POOu1CMuI4NgUi/EGjOCrzuUs+t+aFCmeC4OtIIhnbckgBQn/gVlDqkdVmy7JG36U2Jq2
uGivTtumuTFniFeWPmJzHbU8dtmX2730RCSGnvvrYPYFpFZpEKAPA71BJCp98Z6Od5zR6EwrezaI
HGiZaIWzt/EYSMlBWjj4ZE+eM6iYxpVj0qCiZgqF1FyJ8n6Y8HQGEDcwH0t/WM4/lBrKpZ7C6dQp
rIbkbtlwrMTpNCSPprzNCxLyq3RCcgOuumHwMfGp35Oi7/FgBfvtAOrcrGcoXOQmLkd3Q698OkNI
mangim34Lr/nZGIqR2vGi6rXLrXYvX5vjAUhVzeR1VcR5QSN/oCGP8kzxtPFt0QvoT6atiGgAdeY
gHmkwKHr6cHA6v+VfyD5WnKWyFwaWcl2APfpeQeG6oYsFoxS4mLiMI5S+N05t4NkreZI4bK7kG8q
33TBqPWX8fvSvln/aZR/+PWSsD+sbz9vE8ObyXJ8Yw4r/5VQbQxLM5W04JHp37xGhWQJMUBR7kXg
kN8zW3jhuhNp9Hiq69d0Rv7o+8rQnCUChqGCzW0V/dAyNXCQoR4FXNW5jbShiZlJTY9V2EYWgJJM
sjXzM1rn1AEOBvVLl/mraAFBl/fERSvPNu+MXe6lchzeYprkZhFsTxrGbXN89DIvWo8/HpIA88Or
LLr/lBD488RleZv+MJNTOYchEbwVac3LC0h6QbkkkTTRtATaBCZ10oVQz+sKv1u2M4+YIh1rztJG
WK+qMftD3L+AKJHYFPlARCCzDw45HTffm7MCAZFbppty7eucIocTtQZJEFvrK8Jwonqmw5EjMhzI
s8oNJxPqAUR7GHt+SIA/fWqvPTv+Es3xMvbGEt30HJbo+T/kqhkJTH66SOdvClTJR35mO03UJD6a
kXt9EI9dJkUq8x1aL6T1pGSis+U7iHvqlZ3/bTD83ncajSC27LyXYpTVLFszHmqKsfeT9QkPJYwD
9EXwwELOXDawqYOsPsSaRKrDm4ptKDV2kOCj9QGARxso89oCtLABPiSogVGhiU7QHU6jR0zmFDiJ
Wcr+9Plzc4R8jIRusx0ch6tCCdl4ObELZEBtw1X53UZJJgfwdpaql89XLz3oArs8xrcRB3RNaMHu
w7dWL3lsIXN7o2XhA7BZTkTnou5NWlCds+ESXuoVsoBw9bYdSDvb6Apkb+NvKugXof3IgDBVPBc3
hNi+E9e4dxyv/su1V3rrCmNua3OGFZA2F7O2Fz31xUc9l10Z1qBv75NxkkyqJj8KVnAQmK8bgdrn
YrvIMvK5kWqNq27OI9ATnO7b9hDCDIZWQObSTxk1PKEgoSysbDqvE5Cu5lfE4BM7C/BC9NY1v/eL
vhs4SIFYW12AsjyF1BbBee4ACKet5meyikLsb54A3yS8HDGrB6vi3rfytoSJXWxU8/vX8/GDaszW
hq8YpqyNvNlYTxwFEoFm5GBMeUeaLeRukolDCl+lzQL4txRWz6O2d7NvQdsHRremcEb4vhQBFK00
lrWpvacsspego8Nl444ve3/Aw5ulsNXyXusK1/e69F08gxRonEj5RchujKgnbV2ML6yq7kWUm53p
F0cjFrVsV+ELJwgCFZjAwcScBx++vXEbnuq9ttvIsa+p0K0UZ6103YdI+TQad5Qe4sTqLlpsMHq2
SijuN9hnfM4VBrRmxfmDUuhfsMworBQrn9HdbIDlVHO/sNoaT/rG0XtTNCWx/c1/lvImo3GLuMmQ
BzFEgRGafRFl7QLXtCNOTa9/I/GngwJIWOfzrAMR6os63nR5u2SM2Nr9bDBbLhBhQqmmYAYlIl4+
ww5OfkYkbdO4wn9xyqr/BNn5maEPUUccCAxUt2kXt251qYZvWRXsdjeJFIvfvhUkAeNTO62LZLrl
0Ayloui9t1Fmp+IMSEZlMsoOFm+FOepd5TEGmGnyFXwNuQPJSFMP9oaBeO4q0kZt37RJpFccHrqX
9KXJZ+t1/0o/ybkYjvxMYJXoURTQx43MGpNGeBrBE3XMw3LfKPNNmb9xMQ21mBV+LQWXWgqaxvKv
XNzzQc1HyZpXItXXsTvvGS+A8XKZIEqeHUF5pIVH61Je0qExIuOFSwEK0VjBg9n9QEgUr0LvoSDS
KKtupOvJrk6McFwILPGus+OECK4RMvKD1TgrnLgWsOVCMjpCD4DSt9FxcIeHsoaGDLSx9/tHuS3d
5w48t8D7RaMBhr4j4/CtYnLjxtu8gYiFuVEfDIZYw80eK0O6edTBnYUN5SqEKRLI9hR8dTwThMxP
aBmbGV/k3iFL6ZSKr7Mz92+f6nNRMvC1rK3ThzyyiYUapkeZz6X/cY/w2x+2x8xuD3M60HuRyyNH
QOoAqeJfSOLwBQRBBLXNQENxS80J6ygWQTP9c3CC8k4y1DiJUfOYKSY1vU+rsAJtKPD8NbVjxl0Z
Vohp67HNNF3f7ksk8eDJqplI4xl68QI5XpMxokc1QwBrJZ3U8AgeNoZcLTm4UVqgqRAZzxxcKIjt
wTweadvBYzHM1fmrk52I09L+M8s7C1hzUanG0AO6CL/5MAaijLXeYhjQQvOAiu9rl/3y69Oa7D7J
hjn6aASt53li2Or7rmKBGgh+QAtlXEEr9H0PMIaCzyDtCSt267dOELdfC+NWwPG7gTsTQ3t299sf
10l7u3HK52+bPzxKvYiBvG3UUZy/ISV0BDqpMJeUzq54Fae6lZnJgbahkHkCN5hzGcIySgEE3t9A
ShtpRhfHMzX3P5gFk1q4Qn+t0Eqy+NeTwztzrwvyzVu6zyMsnmcQpW7a9MqSdW9uQF7bRxgWpXZm
JDtkxLq3cO7sdmCtgMt2I6rs1hZUpHf5Dy4v6kR2ducDiru2W2XX18lvzoL8QEj1ZmpAEnGWRu3i
LoR0YQy+iks8LgsCSWzo9DPHJ7WlFdZr+ow6wnsw6D/M23KCXSQcsj9RV5e09OZ7nZTa0kW8zi1d
UO45NGMqzpVntPIEcGU2Td7DSXEO/1NEaHZzSi3he1LIH1NVFiXt9wOdFu3GFfafKJHFKbBDT0wk
7L6YWY4Pnk8+VDgOnfj80dHolzpXTfokAGgcBn5jPC+erDbKUXrW7Colt6UZUOy4dJ5PkQC76Ezg
WjtPhxUiHsrZczcGLIEaEveHxAfiA/2JmZBsbqHTbF8ZRTQzjnM50wHGqcZ4DTncUhV7yriSdv2O
E5x+VGbQncB5/975CWxcfyJoNxuyOa4nRt0nDei0ULOv2GgJlmObEfxRErAk6DwswBWfJDKXOES/
oD+4MKtPtmgNfOwxDaSH9C5UAcQBLHi3K6UWTcst8xSLUeA+xrDWGFZK9p/aKiJPGfmEY21huvIv
sQfSMLRXhEIVP5vojalrN8bQbvA9oh+s4TxhqIp0mDr1A4VsUNUOgSuUMfmFkMEsKECvd1ZkvTKa
L3/uopuW0QedxaUKFMAfnScIgeQku3DNNFCOxFKmUsDyHhlFx6vtE44n2Lp/B9oCKMZhB+HgxS8Y
lQaXQI1QEclwvyBOylsjxyzJmEOHGg4Z7Je0GOXLpAwShtEAYl8O6sfAwsURoTVcihZtBRMCC2gO
HAUupRiMvpgJ5LzNlf2TrUhp1/ydaS1AbVqqkPTZW7XR62yqKdxmIt11GPdeYTBais7NlC4QWqMm
bFySx8Jwy99c6OJrJahgvdl0+PMjQrCLK35mO+oFPe5sRGTNPMprErkTbws8RNak8ev2oXHW4n2+
UlZ79U4jAnVRFi4NY61MjyjhvTL82cZHyGxFiJVD9BmJpS+9x4+mE+T312fBg+qvpQZ7YkLD9gD+
ow/ylEK2NXUMInnn2401JLNlE8osN12LgQ1xqLpX6k7zVUPknibi0WiSot6UG81APo0nYbWFwOQE
HuuWSS11QjRHfEnZMqGjeqKMrPDuLEqpPoH3wWLG+nDABmxxyKHuQ2xygwhuAj5q9Y3+6c91G0NC
+z3XEbM/7qSe2dNaA6kQN5hU9J1H6QuUUOggOFqE/XtCvBP9xiDGN6QbQiFHZ1FpWbEPdBxZpALY
aAlk6rU7jF6Kyi4/MlPeVQZOG7CYyuXPGky0SaW9inzEaKagvB0yZYei48H7EnVqfjw7VlVpY2Vj
xu0Y5Qid/MpRp/LYz230RC5kkLRnmTG9uUcd2+R9T9IztwUzg1e0BYYwuKtbbQdPUEGjuEeFxrGa
Gn1qw0oKa28tV4RP86YhVB8QyKi98mk2J6MDQ7O1WX7IzqVF8469TKlsiy4CDM11Ph5bM7NFuwEq
GSHjTkBBsUzCnCiql6pWqqaXgjWKbLBshFu3BtYUsTS7JA7F+aX/mqN7MMPyM87sN9PmBfNP7i0G
OROD3ecOHj+fdewZvaL+kdPDVP4hOWMbPT+zb9phRiPcOMh4x3lgBTZ6IcLP2jnBBOmu+vnzXBCd
zOg8MUSvRI1hDyAeX09j0i83KZJYMNOqyV4C/loLzWHWYDmtZHDZhk6Vd74CkEcn/iAAmBV5zUd/
bPypDqX9rc/laZvQE1VY/dT9fZ9T/MhlVDtuQEBGxTZ1wGhqq7L8CGyUpBZMgfWXYquT7o4rMzLt
VV+XXxM1enLIdXR52ZxREeCFvfxNmUCNG+RXpKCgSsI+DSvSfX3xlT60MsF0gbpigvZibq0w5kvY
5uSGrt56pSrh1zypvleHcMNCVrFfXohjDRoCZ28Qe6hpZtojuiH7GRhJ6aM7TQF9P93E7N0nECSf
Q5FXCD1AesQapb6Eg4hfHXDpw0Rw+ycUAlIUbBTSVNTe1XvFKaeWu1pQfx8HhNBKKT1UESSSu576
zFT+FW1z5133bmRe9hdfvBr1qywHrNnYGJhDTboavac75DOgNgkKi5DNWhal63Kil6O0ZfCMdOry
l28wjTaueznfOm1nhd6KKRb22b1GDMfU687Mstc2AHmMZoglMGgWk/9aT2pusvXyIGHA3tP0CCWe
CCc2Xdbd+W1AFKlPTKf7yWT3Jdpgs9vPfQAXtEycEQjw+R10LR2uJr0xIwYK1kl3B/shhX/H+OUS
OIbfZPGhLsWccrC/42I+honCHBuwYbyDOVDo+SfGDehOK2sPQiB+SqhyYEDyh27m8TbFe4RZrtsy
wK2yGWMhBm3QmxuZhDO3TF0FY6u5sms6Y0oOlTkSD9s3Aa+WMm0BAJKNtjvblWJz75IgeYjFgM19
o2QIq8gAo1JbuaWRVDbFwsklIhBWiqtcSWGLuIF/nu0cbTjFigkwrI5whWseZJ04R9M90S9GYQdl
C1s0Lr6JaLNfoDpGmA+HSj/VGuau9WdsSqDhv6C1h7IPR2G+5AsqEDIJRyQ9Zbibx/Fekpzl+oGa
CZRrHVJjMWWXZTTlRincxnNrMtZ6/Mlqsfk+7Hx9cHFlxr3SQchbOEQV/VvZB++OaOhV49xjoch0
B4YTbHPPZ2enZv4ZNjQk5lLfOwLEczReSuu/VFzMedmxBG1QNRbrDNo7nJdc7uQxb0Jgu/owBiIe
vXSAS/xGn71aqdoAS3fwHrAecqAZIZFIihYyhDJSIGC1chC3dEQem6LFNBOe4K6wtU3lvO7hUHHi
DrlFTaUeaGxiWNxjlUjHJvb+OHL4SRgxm1VlbRCkIlF7EcigyclDLNLqU4LeWEy7BiHpoCyX7OD1
q+zh0A5y/B9ims2kFj0vvOUS/SbirAc1b3lGx0zVUQTJyGGB2Z98lmlnzgb+RP+ReQrRNpWYklDu
tdxJIG/tV7zAX/LvRWrD2VFTyLyxuuN99evfoOXBGzgb72MC31eGtb37QSVIFGL5r5YtK8172uhm
NYxFDhsDy2vXfX1GQFyKPQXIRYVD1HWsdyDoH8hXWsB8RlY2f0OJvMSYUUUh+FqxY+UZzP4gxvhv
7S8OZC99Zf9Izwh6+qHFmlOn8af2FQP805FZe8pVQVN1KPv4BZieDKim7vM122l4bkNSBlm/qvX9
Ag9cGaxVk73NK3A08DWuSuoiiArK9ywAa9z7LMeQHEx0okQth2O8k7PFruGc1SiyTStJyrtq02Vm
NsT1VSM9ApRg75auKIU9FrfGQag2oNHAHm1rOGjJ/+MYvFIexz85/bMllC/lgZ3i9zA8I7aEY0H2
ULla33UIu0IGp2gi9TsQSUtRVyCo7aNf5yIECLO1cruUK47hjaUp7yikcd7mdtdxQgMFDByyQwfo
FUfBOR8/k8wKkMMkMgwaQiQiPIbaS3kgmPWBtkKenZslSIkogK2gihQt+/viYSsuOU6jd//lFOS3
4ZF4/Iko7dRYIK1mXTFQr1p/GpfImcEWx4w4YmmpqplLR2iCTrdIr7Cm8724WKqVo3yPCM97YDYe
nHxebIvPfmA1iyAmRynGTenOcIRLPbFu5YLsSNiBt9UeePXxpjVfm+deHI5LZmlFhCFTdv8iiSDz
EnyYjrgEkD9uNq2Lp7iMcOk6Hy4vXsrK+EF+V3pcxWsmcI27U6+pqbCjqI2xXZup8q/3JUrNoUC0
U81GbQNKapZwJ+JHu3izkNTUasAoZpe2cXpKNTiMU3s4qHNhaSEtpgmF3oromEgWSnp3iXwXKBt9
uvvfC3idEY06xB+APqm7JzRDogtXeOMi9wrvUjf7HCs/jaMIt3uFEhNSzFCqcLFsEhjjL2KKxYvX
Uriy3g2vO5MXG/BsRrjGwGO/qgAr11GX9zwHxgn5TOF1cMoIapTmNez0W8hpUOAJ6UIJJJUAlzCR
+8EoPmPpSMn3Eyx2tDxo1t68UpxAHVQ6VlZNgeGktq6ZM1eQ1PEr5aIkzt4OLT30cGCio8BWT0kx
ljFDvgvcQOg5mFcsn3FGFHzRE8EBho70tzRpjkZ9KVE7AGV1n2SlKa5NNYbNjTQUIBE6NTM8wDOe
oewkxrvFli2aGq+g+oSuV265QWJVQ9A0fRjm53e3iriyUa7SIEhnKauASdC6L+Llbrlkvkh6l/3H
PNMhwjy8DvuZCIVVNKs1Kp5E4RliyDxgtKl+6VudldB44vek6CYEOo8kglkmbJitKjddjni1OnQd
MIDFO9ekFDyC0wQK57JaYYh7utQAnSMhn2pT/jo/8xvJ4TXdb8uoyfy85MMh8zyqC1NINeWnDmZT
5tQzk/Z/2q984KtxCV8+dcRa5SGWFjHhE86FjQcjrD51piGrRrHoTJGTcqVAjjkNAYxoXzsUbIcB
olUR+jDX9mQd5/u7qvSalkNrKguy0pzXJhl15RthaSmG91PXGl8jQuffJpkbCFfC2AeKXq4iQaEv
Bg4UnW8CJyU4GRVBH7vB/Tt2erP+aJC1CWq/cW3djabXyg/GVdc1vtZfNhQGRXRcIU03IZD54Nlm
ZvBNk+Bss92DoIw9f+oxtDCuAAUJ/L/ej7yrCkSFWfGreGHldnSuePCuLNL64l3+LhCCl/r9qsh8
K3dw7A8VlN2tJN34neVpnEjShejZ6Hc9nMrx7/kv62iTX/4DVN9J2gBBFprBCQtCKTPLmiRLttzB
Pee6gQm4VyMi0JZPiBNrf6nFsftLGcu1e4mLdiF16mhpv1z760GLBpC0ecNQyDtnYxiCq1TOi4MU
lV+YAThd5h1PtCi9AtqLyJmbxMWWwE538ujGGXW++7f+ZxD1g3kVkTzGAA5cILuczIrKpgqZTL5+
1AFWdIHV/6xVY18Gp+LoBvKJruKT+bApkv5+nQfQwj3gPuabAQVF3ZSOgZ+RyI8pLzbAmCaGhEuK
MM1JrUngBxBQg2IkAJ9cr7n975xwmMJRw0xZvnKwDdnkYpPil0fLBXsinOgS3z1OdWJbLmTdR61X
slxo1h51nvCtrBo9iL1tXcroC3RRZneX1qfsidKBxmha6mNyit6Ax0D34CZe5+B0J9qWpaY1vDVp
/9y6Iou8XTdCetn5YQOBSIDV/1BQlu3rTVprv/KndDkRwZ/weBKH21XUFleZXwRtAPOadrx10IcV
s+zBBJW7RksDZi03fkBFHBOpuOTpTTCeBKaI3/hkrTE3SQmP8gjR+pC7a3Crqu6Bwe3Sy9TCEzvY
OK9DZzdBS+amR614VvDzcmAGoqq2Jd2Hj2TT1S952pREQyRhjbbuHcnBZnLBAyzUiCt7eYKJHi8R
kyhXMj88maOCrSBogljPDGVPJHzFm9bJ8tmpJk9A2RZK4Rv6O9YL1NZMhRXS3VifhSMXRRJbwhQy
BGReSjwMtxpOcVYXAslEvj2Z9nBw/Mtso9HXiU4PB1y73ThatkiqJc4QT4ul/o3sHktkTcFjd5KK
OriwJ9xQlkRVzOFBACObR8eMJdgFcOUvJeZBKBqqDW5PYpT5g65HVN37zh4EeM/3yu+jNZPWxzOn
SCFLNtvXNOdIG+4eb9vBGVIMQS6RJdIjEic9fgkWIDx0HjsRLmYgEiDg9VW7LDyro2nc155Z3/8t
wpjgwTWx6sctbSNiYXg9KFAS2knmMStkuKhKKNbJGv1/53J4P9QYlKgUECiZ+H4zknWdG3hCePfw
VFTZt+DyjV7Qoe0r5MbyEBsfcCMEnhJd6UpnA3wuPsoAuiPYfSz1VRrbSAw7LfsMlYEdyfMFMpE0
Eb3WgJbKVjptsX3hlylT82fINuyDPQU/X6bXCZkDuYH2CbTiXi0ImnT833vZsLlFhDf7imCLtOY1
wQsk/kzKEA1VgZcWI/kvd0H/Txz6c2radEv596CQjuCIZ8hbGsfa0R3oAtlbIHluSiY9fDwt1xN1
9PfIAw1lQiav/6vYHl9/XdKwnq4Nw/6abxr1K9xXT6c74slvuwkyZxBSX91y9TRcIb/CzzY7cQ1Q
zKDeHw2Jp21T816EhFhSs1Oh7guVy+iKdrhrL9pLPa0aWIyvh5vEwvhWbj8NsnWlR7pEUuNAGOhb
A2dT3nhCGNMXgyMaRGfEDfKzM0KHwFDUMFFPIjmiU9QkgzctzkLJg1T6UcOUjIFHBnK1pLKjRvd/
5BErUHByCrGw6Kv4uBu0ataxDrRMsumxLNpiYsS1aFzoijhNJs7K4212+WcrjwPJ5pVr4urSKzoi
NJZg4ue/fmZKR0Vft11/4qFienJQZHGNPDowHnY/kIQL26EWyOGwGPsCIHgwm0RC/CPXpBUoSJvi
vCQtbgNUjGQPlFbKZAl/aLCQqJSF4vHrzHW+50Kc6Yxna7WfjNE0OPwIsUjVWl9H/6uj4Za1NOES
v/QZDUR0D8+AiBM1p94pYrL81haRqQDVnus8G1/J9lUggj+c6ZN8lJ6il7HrmNCw3Lt3aF5Qo58b
sNAgJ2m+CIck7CzpPRXBCAKWrfSpZzyIzk3UnKVm9l3jzGeFzzLHpJDkh5QUAjsCZwpQlMO4UgqU
K/HGdXqC27Jbc2JI8ujNeEV7mRDKzkW3+f30mhTiKGD2/ts3NnsoTGtS78PukvOYZHoKIFQlr2G4
LBjayxuA7m2o3oPebSHsPIlsYRM2ihxYW6WE0wQXaiDNrtwtTejp1RtUX3g7g+9XEC5B8ccVPW4i
2KSPobvQ1DL7TfjljsUBnkK97JjH0nKYGMCbiuHaxlQqtXEDX3IWoA1qZ6dEf8g1ZMbqU3tWCo9F
79YHJX2TukWzvtpv7389mFmgVOTl11s44lKPoh/43j31Xh8brZ8d4AHHe1LFAHarxa/W+8cS1b5a
BsOXVtrWc3BxP4KgxuCwwi2jKeioSqe70echdeTEvIiK5Pxx/123D4eA7HhIOFcrhFVJU/2WdTf1
IhF38yixtFPxluC0E9J3uz8jWqT7aIHuN0kJ7xvPB33Su2xAIRjXpzbSZTWKLC47569MhwGdilIe
u9cjz5SeYTgENeXwH+XWIimi0m9ixq3mwAMKMwf1KSzLP7AeMXd3PwgKvpgygCsIMMuxuewHYv+K
qybxk+fD+jcAuFMxDDC6zIXqW1fjGFV+aXUcSnjdYHYb/3K6I8d7Lo0DMzTW0feZmZQ92ATgR4YT
GyDGAeQcFXUHd+Nxw8y/39O4XLumJJLwJdBZ5edoSJTKogeUHj8Anh6kVhtlkU0sPxBUuJa4EJzK
tFypBc83mPezhtPpqseH0mFEd5BAkuQBgsfJNgihMTxLXJM00AvG2rp5GYdTGwUD78WBFoYxb/MK
V4b/VxgjaRIrL782Yjb88HYZTDj1JNDww4HAhspW1LIxInmtarJsUsN5eKGb3x+Yi9AYcfyH1mDV
6ITuLHNikWs+5m/l/oxvHhz7DQwtbpDJLaQcdVyMRKS5a0T+YRF+YmhK60rdcbNv9DTIFJWdheV1
cVhMOmFcTbSbjMaIo4PxHFXjYMUwt5eacKmbNgNGBApp1uv0oSH7INl+z8TZqPxXBv3Jwl85fVCj
T0vkwKIfCfzpWEb+QNLAv3SPLLqoPKMHN4zVfNgm8OjelBUbTL4+FVZscn010H047KjdMGB5tM5G
swA25j55SlsKXJjrh3WnLNKcUsPBKnD0VZMk0pgsI9NeIEY7LkX6/jv+45RVi+XefdQM5ALrh4/e
ykyYGApnJ80U39Dsq6lfhOHcuqaSgdPq0A+fDXOMCiCVqLWqam604KVi5+3Ysq8GK4Gbk9ZVxmBS
wtV4ddBWxhwLQVhqQD4kv5VAVaEpLD51+I2eX2FbAboWwkUzLagRoaLUlJZ+Wfhzijmh2UTAXywy
K1lKdsNIJpFmIhoABvrgjewXX+FAiFqnKCnTbeCzownTBp381xH4DlJlt5TPNN9XxyHPRPoBw4DF
Vtfn/T47fM64U1Bsr9Aq7h/nPhPjWcRkeWsaL1QDNniJ1tHz/iO5wb1bSoG0DYKdb0DkE7oMI5ah
MdZUp6rk4JVy/QETJyH3h28jBOuHVvnueVS3j8MdT2aNHj+OGKbPGY69ERlv+vi/ascQEUFH4dSi
l5Fqo0fLIyySHXuE99jRNFkbr33Ho1AvxbgWzkBskf43csnTXaCk8DUNwJsoshLcgEevNe+XAq41
TIjkPqbZvSWsNhkzH4+VzpVH4CWgq9yrZ5HBLEP1Jc5qJq65m/9V9Egs7xDOzVtWQd+osVQ6lZ3s
UOyVeLuqFG/6BHpyRqO+WPbf/4ZqbnyMkGClhJanTEZiNEAHAwSdxeS8Iu6YYyH34GQa95Pu/j5l
FF6fwjcmXGoL8cURA2hM/rXExKFmSy8K94a4QN9PYfw+9lgHgqJdtFsqgJ7T7Lb5j85/fIyCATvI
YveJZ4xFKN/2oLnTq08KLpaFZNJZh6saL/xktr0ek5i0SVyhWtzcWGm9zcdhEOKgKor87V8A+i2x
fkxVd/+ekZeI+n1qcqHNYxQEAHuFXL3swC8Wx/MAbLCIg2lMAUjdo3lfCk4JLtyj/ZHUVb3H+J5/
8ocWZkjXKEwbHggiS5aQK/LGnanUVPq7qKjrcbDyTYcgBKj8f/Fj3vHiZ29eOkuKCLXAHhVweZxa
xgnjoNTg8X7VD+ogcx//fRZBOLcPbSUceB6VFHeh4BcSrRwkQVpJy8zTWySEmP2jAU714Lar1BMD
mE0uSDnI5Ujkx0ewZR2nMWBOQZxUUma0gzXojmebjQTeeb3fpgviB0jPvxHpjfGOPiT4kC3LKBKa
Fr5tgBcPXqCsw1U+OVI0W9oyBAG1kI5lZQV3LWqwQbDUBoY/oIDMOX3ikcjY2MmwqZDVN22fuEh4
LuFEB7SBdxQAjmC1vScxUfYrkCUpXX8GQ2EPCF9M6di9iWJyS9Kpnj6Jju2Os1doeZYVgMYkI6FX
c7QEjnPvZCSWKgiB8pvteaZyi4owp8RYFHiP7c5yx8pkHp5BQIZI3CSLZwXoBFAh5c2D/JD+EHR3
GxM9l2vsxt5lz7wkoyYJo4lfrwAwFPQMcXAQofbjw4fwGh/ms6tdTTnb3YUe370g1CBoE5SgMqg7
2BIkerJTp0sNNLXY0BVZJDRLL4hnll1dT7EmBjPB5tNdEsBP6RSmJsdm2UC5ebJIfgRMxeDDPYbW
FO/Tlv4WJqogm7hM/4/gJMk1jJk8r7KtERPKAHc5QJfmEkwlY/VmMDA1oWE61PzB8iDkgP0KJmyz
+PmgY1SUDoDKWl637sCiHdBtNzP9uycCEkURGmQnLQXkOmYqXsR4mPByrVh/uzAcJeDd0/SrtPXB
cQM5VyT4X0G45i7zFw6pLWcO7kLGDVt77CmyWrzb7XBetmoSiDZLtDQSBwLNL0h7Yg7oORbITiAO
C1QJBVYgilwpSZ6MoWD0Cs5//08ukpjLaM4isM2+7VDqyLnqQHRQV/U9MfqWqRu88Yr276sv4bli
LSe0TW0R5C+WjEedA5LinKDxBVshPX+m3FxKwQu+oeOORYw0fp+jCTviZrmVDBLOK6w+/1iLqhy0
rPUCpn7YReJk0Uxwc/5RZo9BkibYORk31S/a3MVDNLSLeTMsuECloi9SbjSurdDm5BVBymUdfniR
V1r/XJqXp7jywNlalIYw+Sn20GwriPaVDzrTGrvRlpwXd1L5EjNOrhHBOjhQKz4DHUBjwgZo8nt7
Qj/5JGabE9IQ1vygpuMC/5YsfClgMVCdsHIS/zpstk2dYRLI5jODRi/AHNKMLUFiXGSI/jczwNRA
JqGWwnd3mVvW6dju1xgCeJ0T0GaXu45aRMAmNci92sLTR9qWsXDSuBLfevYQaz0JffkBELMz+EZz
/jZF+nW1gLwXVCTM+0ie4khahOcXDKXhxr/BwU3+VyoVA0+cUlXkn0Za8MAjNItPduvRJYbdqDqU
WvAvo3ZByRg3STNjWWXloXoX7q6J3gi3rbtB/PTUMSUtrlhXo1Fe+dS7+d/s7OeN3QBEhPLwXMDJ
t3HgEmax6/EXjRINld3M0mqIANSYPe31e0/8LrGBuFoCi6svhwd4Reun7ixD/h8pAoY5iAj4W9wz
1xuk4XisTtDVc1HkJ/ubqquk9hSGmsbIsfPotcK4T33dpcKp+yKKtMOJesqrF7TV0A1B4eV50QP6
I5ZAeRsG5EoWt4QCxFFPUPgGjl2IFQRkqQxxHbEclGWaU809inp/eVXt33NzWLaP4HbnYLzJEhRU
qX1PSjeBpDInFthQFVLPRvDp9jFYlGMuUkdSGsPzmmyLZt8AfvzJ9NULQ1zwqJNAd6K/j9yEi+7N
UknpCJ6TFMU2D+za8/1M5gv4gWLM1izyFgqpV5y8nOLVHuECrP+ixdJBaHa8Aqy0e60KhV6LVdQn
xrBBBTtPhrYVL6Prdf+LiKRP7t5e1qgnPYG8eDDBzPXwpS2+6xdibAM/YETXS3WMZlpxh0vcUz2E
ZlCUEfCPUfh0Da1HyF27/YxPgYsMEw7G/OX8FCnBO5Hgt/Tp742Ws0IS0TcZVLdarfHwj9x2zuvj
SVWX6Z3HmoBRLqWyVbr0SpPxdX13kizWKsQ7MrPuJ4uEW9wnVqnuEi057hDHTWUfNg4xZqewKD//
3eYS4v50l09k669W1GIsOpAQU4YxrNw9dqo/KEJeEsPllsNVwBPM6Hy1nDNmLrHH2vu4P+ZBOheK
ZJCNH7b+tngVFIu14yrQw7woH/+6qaGW/c7O54V4+mxcGqD4fDioUKbjQ7lsCD3yKCHfD/E8ZEwR
g2ar56GtLvDSIT5bFfIGJ6HaLk5ePLm7wMnH1rt6cLxOD/i1owRwvM0+y1BlmGt03LtJClZWRWXD
BdKzBtBf6IU37OxQABDwceqWwhIxEtYMIdwtdVS34SRebvdOrBd4u0+YpWebd055FZ7TcVXZ6+xD
JawIyZm70p9qSjeOLtruddWv9g2s7VxXKj7jsFh/pmjnSTBief7GI9nTo1rZjUcRZCdgENbtMmEC
Org657Su+XZKjmrL+OICePROJDWTXbR9wFdiajeiLoJ4qq7YhPOE7YqX7NjsmrSngWtEvhkffcAF
VylFGG3RcWIbQ7dm4S5FKAI0NhIk1x344bmAxI2t2gzkQYacXx/2Y1mtJwqrUhWCc01z/oOr6O9y
J+FBeQ3hXM5G5UsEbfBSRfn9+RZlzwWRPG1ZBS52PzNoNtmMk+iANKqMZmuliMFB8QfusN4KEt9U
XxAwSIuMDMhiquv725Ms3kWyQFyT9JDOD4WDWXqvjzNDOS7h1oceurObrYLI0DxxwaQaTgH7kf7O
veCTFwn1DVdUfmRPrY44xonIoPp7Icwosp59PadKuuV/TpSFWnzC1H+shPJ6V7NoWL7RGuBA1UnL
wXIxF1g2MDhExwpGk9lple+5CEUxc18IunBCj/7oS1VOqXXYmZU4r6SLzK/dmphMpXtdSEqV14ZC
gaKFAIrATuVkmN6uv0eHAjhPytc+sb+zkfi+ODr8guaaqciIj7DOOgc2gDSU30tNH/BmlijN8Znz
iAyWmJ2WtljMTXdKqSOa/jpytfoMT+982bF4xm+88VP6cp/u5Z91LEqwUSeUMIx4DlMwsdOAdQrX
rlvP2AiCyQvjhON/EV9vgT0EX/jO22PHNIS4rFAoeFFbwrNVfdRKFgpQRUh5RDMZ/xBdwBUEY0/9
FaKI21NryFZoMTpEu8BNGsYrnJkyFdAZjxdwCr4G85nt8pdT2gCs6qr2q+fx2/Gajv9cZsZcoUDF
s+xSKJiD2M3VpyiyIaTCJCv55vNJoG7PesolvP24tML6+9xOEnXPDR7xyud3K5fMUvInyWRJ9MVg
AOQAVRvXuQa7AimEiipEN0n70Vbvhs42kX5NpsMRmp4SyT5Essd2HRIqK0w11Jkxppq3QetJVu7A
PyXhEYdQ2MhAcWF04OAlYG7bNpgvmD0F4UGkkWyQxbkOYsfDRuCSmB8DVxjWG2PfijNMh8KCAYG1
etEe5V3TJ2YRGhCwicL8bivjBV1x7wbcdzeqMB/iVocDYAYy5caq2eemj+rZzgcxTRkghRU7K8FQ
eqrk/Zkjyx90gQGJxVeIgnQX2jwx803ULgPN/Rtss9fRtd0RiB9ppcwyMviSnX9Y6Vd30NiPaIrY
xC2kH7mu2QUlUc7oDCEoZTtRenrwP48/s9wDgJRBwMfWfs4kjfTYuyQxTBKjmfK+mZJzmW+upuwz
LxLdWTwr530emjaOEXL6raWHJptlGnDdiOQfJZ9R+1r5pgbQE5h0ZwnZ/t+WmdwfDAMP/B891KTY
kPOyS+R1WOyAUZuPyQB2ZMaIBQed0UWcDraWbWP0weHDqMhyu9IWUCXf2vtQkV+V4y0kX81NOraY
SM2jWykPlBAYqZIFyUOPL6VvCeHwp0oco89zsCoxRqL9OUbJueN+/3nC0qe0e63E2qeva3U1fvTc
OmLaRx988BWp+5vnwFYuRc17W/vrmaYhrP33bTgdA13iGvbnshCJp4Z1ijVQ9mdpZ8v84b6oB0gY
7rgWT5RUMoNYQcNxRlAd/q25M1KJ+G1dyG3YvFigz4RNWU/hhHV5FamvfXAV4NHaFkzUnrIMIFqk
CHiRlyVQU3lgqq1xQLwHQhfkfqVeOL4EpoyCFry5+ei+S28jPcQTNHWORWeaJZd2lTtTvPXX/U9k
Pfa7Feifaf4CbAXjPnWcNcTLA931S5zpXDLBlsEVswzH2AmZ4fvbQF8ko9Zg/a0/Qr97tyUj1YJl
Yrw5ERzdsvv/xgRM3Mam32yPltUtEzHnx8rB47bj6Wfupqd7k28+DbUZJWcrmGmkAmVWYhlBIepv
SJ1fITF14VBbWFip5/EWk3TJUjjObkUKfCVDC2ZduvZC9rRccss1fd/1LBvuUcbKZBMC0jiyfyvO
YSa62oJbVoO6Ig5ffXf3BHetZC4+kswbRaAntpVhEts1pz0yxXsp/PrpuqcLZeX7r3NPVvLE8CB/
20gEgZnCkFeHTmfNb864AVoTIlP82GF8youTlA+L+tjQTA5h2xXze1+HpAViB7N1+C4OMqIi98YX
9Seh/jK0xHltzNXyrd1eH4ZRQWXtULOiWoO9wAhUEAOfiOM92L8gKEJqBBD5ykixzb3iLIIF/G7r
DYoWBHOuyS5+kn7446si6dKgA0ibn9QVA2PsrJaF+aAdk5pMSDDBfFp7ggNH7Fy5sgZEDFF6gSoy
1WTiISG9w4jrnmtJTTWkMyf2NlhktfL7FSvRcmyhxWgkBC8EvcteTEyA+IopW/R+HvErd4Q3Awkm
Zq+K11GPv0WJchU+3iSNMpcyIbMLOcezsB05ntMWHO303WfDy5Y3eBUVdrG4f4vndUC1NJAP0XVO
eYBYeMPJLy3RH9jE4rG1ADHYpnAZdGUgqchxs+J7iCRel9qGMmctop9DGZTctXntL5tborYIyxaQ
pLBfERPEkUwT1PUtrFpX00zZZ15iWjb/IAuBeUPY4MU8uWPI7N04Qi8sZiTJZFOTJ5Tl8Y3qF7DR
jwxWUX3airGDWIdPBR41ngriLUjtug/ivU7CjrgMXh56EDJAFsv9RjN2xh7npHr8Lhnl3s+hSgIS
1Amd0lyGz7ArVSblfwbIjdatCQt4KMcaLWUm3FT5CyWj5Ei/kc2ZiY/GpWPaWCkL2NbOuf563qg0
C8onQEgV4eXEY83a0PHA7XOW4y68ysfgwBafOKvng2pHF3y0QGG7ZsRkb1afNiwv20MZqNevSDEh
K5zOgJOO+eHBjeWI/0Dheuqe+Bpna+MYIpCogndPyUIhlb+dh97kkrLQ8+roAMf8BPYW/r4D3jAM
5o/OlbpO9ckuLpZ8FPxQsjwM6cfdexr23bh6SCYX7H9D1GauF5tuTIVpbn9U9vjDAaCz1KF97OjS
SgcU6VqtK4JAv86/PF+jZWOjlFHN7MzOZf/LPSa+L3GfqrGkcrj13FIMMee5HOeIwU5Gii3LE897
3B+gwsBkoQi3mIeLk3goOSvpafzdTPX8NXWUZEOiUNl3RMwUp4WXQfwH/aOfeYggzYkB0TrLcwRO
Biv1RXqo5UWB/QvpWSzYwTYCodr4m8AGrM/I8MM2XzGS6S7K7sIBcE/FE7D9yy2q0b+zKQK05hFY
VCkp8HT1oNApMJjloDZR3+9hZjAPad1vV+wu2M7NoQ+FrnYBNNAfal/efgzba3P/rHsiV/lUvC2D
Dx7J9rhGfAlFUk2BHmzFyuAEADxa3U2tksQ1hnKu7C+xt8Gko7JsIsGXiWJi3Nt6cyUNIF2OXkKF
RZltpdkn6gMY3T2qvCLCZ5cdvpz4RH9PuQE+Ycs6lv4eU4jPbTthbaZWzQfamjZMPxPvb6sQwD5U
zwPEyHoIqhYU/s/2TJDZAWgwAxcKx9NMhtowhg9OooAs7mX9nk80JkhDySMRyJEwY5fuWNd/8EKQ
FJTfqtFF95TEUBuIDeQqaK8StYnS41jwhlFJQvx38Jb34vPygHS2ZmfOP6nap1x/sw0Vj13AiMJJ
1OatmMaoXRhaQ96aIwsMlFFIw0INGdcRGc7T5EmqZ6+YVzRgnKZsDIgBYAGq+kJ0yAABqYkvb6Jh
xdjlf9fezvnJEiRH63dMwz3yFATjoGmWkOWdZrKeUU4jN+NLYmuf0iefPd58qCgtDepa3K2T6LyQ
G2G+Q7t/i9ho8Lt9/cfeD7NPBgVqIyp6BXoSprIrBWLSVOtspIXn/NPoNQSEPSz5ZGSrSHEYmZIb
Cmxc02nAiS4BFSHsaPI6WVIn6RY1fa4sSHCxGgbPRrTY3KxYqKmx0kyJ9qXdAVVqWNS8ZZDcs4ZS
M/UX6NksU58qP/B9Q1K+NFMxA9i8KI6SCHmP7UBFUz2YsE/N2QR4hoK5Gbr8xCKLZ5Y5k6L2Sisi
bGdOSTVAFcwK86U3A3EwtpICaREMuj+hQhz2U4sSXgtijsOU/dG3P004CTVfFdz6iZELzMwZc53U
Ss/sOoDr62yJ0UnDbR/7qENJvs/V3Z9ehyqvsdsWLpZoc7tjLTFBpseXMPkcFhjCgUs+sXgUUJnG
9Ri65oBgEI/GxhmTvTgyZSG4hyDfWLVrwUmryjgw9SSt7tFZ+GDZwqY5UKFd2fH2TOn03K3gOCGx
vhlIKgCdBZwyQd93cFuF2ixEDbisXHsg57u93zNrOisqVI4ka2wwlW1yO3gLmf90FpXEhfO0AWS1
/pA6SQIrgA2FIyfa3N1GGjE4LU40MUD7sK1pgw4dP5QY0aZ+Ri5b78WuhvhO04SqzIMbgrrcfCJ/
AUV5J8ZA5wftnZF8N54zXkOHXQwWCIGIx12SMjNIwAAogGR6jyoqnAZheelCjnp3x7DlMEjcTVM6
rmy0ewvWI/uFOoAr+XyX7mv7Qzld0fmXdBh6mL7/v7MUn2N73L9FfVVBqaKOtyYtngHktf9oJrNB
CGLolPSyy6QUvsPkyIvKkoCc1Gnwsg/4pL1tOiNaxLk2dg8Mag33r6SfONgzkV8xZS6WpNz/YXqf
cpvT8pC+rwlhP8BuijWjKjVdFX7PEQxQqlWeXcH0RENoUvqm75ZLBZmL8pJECkzPVFbs1kLjFHsB
/oqATE4zEhAiSu1oqHD5IsKQxIwBEISBnMzcdVi3BWdNuRkiIiHuZtzo5k0wfw5D2b5OO/fdLfr9
3EGGaayWbvL3Szkf1tUredO1aLP3agl61SCcNxnBTyUKiIryujli5mncoO8M1u304cc6oPxarfsn
2/VehwaWxiUp58PmVdKJB9d17aZMGONfjY5tymGg2VnrjthAIJI7w04e5Rff4QwJvZREC2lsG7j1
E2xwpgFL+wt6bvQuJFpwzR3vpyDg6Q8HkX0EsZlf/5Dr0KkbiZIS3TWSoxMPrqVU0E6i2DchVaZo
va7FjMUcUOOmrcipCk6E3ZoaLtgS4MMbZNOQXE0/f9G3+4ZP9ponTF2brK4jI4Xg4122f+8xoOxF
my6OTvwtdeK9e25wS4U9Zvk1Hfj3bnW7kmbRjCA2Z/ssmWG7HpWwpD+2RaPayiCxjyAJYxV/zJ6R
Kep9m8mosDOj0r6QcDa+vRsrg/ZuzDWblDkBRkGKEpVv6/TKWFRUC6nu2RQG0VlT8c4ALNJbasZy
O3N8XznoYVPXl4K3qdweTTAgD1ESMrtq16KSB9mZ8yvih+4wa0ARRNBjXwqRrnLaTJS61w/O3iNA
ImkaYb1VY1P3O1SroYKFJWdvgLsUnhZLzDxoi40ypzzQfbNkjnxKPnog+cYU72qmmUfW00+WnLGP
+eKewP/kUD+VcOyn4Me05np+jd/3grugWB/YrfEPpiGHPpr7zTcqwjOSlVruDNfpv9/Q4s4j1Z7A
VJYHcayamQNXTyM014UXmRW2qpTsSWDXXHxhFJsrfpqJhBjP1VsC6MeSZs3fYDNJYrwrK/ixnXE2
hynlkjtwudSKErE0+m452hs7vjjZEagB876Otzgtxa5p4u2JRCqZ5P1rjH2jXPt2v75B6SGMHqVs
T2qOLRodJOtXRS62Chz/HwfarRdParQ9C1yhjAPPuYtR1s5BDf62CU7+ATE0/iWOOciMHars3BVU
wzwsEBh3FpqNcMDavWHhYCSRd0AGC1gCPtCh1QZI+pPWSH2AZE1CYb/RIl+BgLzlv5NpDKdoYQw5
nsv2sbSud4PwaKghUBK3Oe9nQdCz4cESY1ddrWThSxSq2/XLYgQX1xnMzKNWdBD5SorbLvbfw5jI
RSlVP2bAx7cYXb5399hbCBlkgHlWTSfT0jULaK+06tOuYysBelJWR/wY8jHfoXD7TM8Vvaf51Sp8
7EvZpp+luX6Tqir+M+05VXdnfu8ESCvXm1T2erSo9ybHmw1CqvH3AplM8pX8iwAbbDWnMilJDsV4
QcZJE6rjCaX83iKh24/zX9EL+HjEQ0uyM+UCezY/fFy5kyW7VBpzfpESqgeMN3hXIojTlN4gEVSK
Ni/CvnV6Jp+TEL9vKK5aFd4DuId7Y4uDUVx8lqS/IHP7aveNe80wZqDHj9PGXgS4vf8N4RqJ2KfO
V6Y7cfRmaeqy7GoKk92dhplWdzlhzwiNJmQ4FgjJHoiAT92kmgDPFxJbuFokIo6lKDRYTRIR5qFz
y5dcUulgKm/VvahLYd7D+UYMbKv6ggr+uPuHMU14j7C4IRCR0/GSAXtgFRpsP3KAdyABMBdjiqEJ
o2ujHLA0uYLJFuQJRa+JrKIc6o6phLH635LIFXbDsi6+k8SGEmWSNz7NLmKGo7d5rD8Nn5zyA9rM
Fr5QBHbbmX/2dNbJPPmHFiu8F2CV/jiaAlPRbEQXe+7UD1A4AVhxOhvELj1lWY7OUSHgMCiplZuf
XpzTWwHFUXj9phBM41gSEyJebgLZMik5mhm7xt/MwUOgy2mhY4EEIoyKfUUpDuTk3Poba8vmKWh2
LdcdHFlkT4+R1M3wT1QQtENOVXWdF/tzuOh7sq6tPu/DkKqp98Ac7t86Mp+DlfI8NYuE3BhGbjK9
FOUYsDvCI3frXxmxYgB9cKD651ZEkCEpTQP6W9m47zVB+hEldDL9xefal82H2i5w6Dzel5O7w3DV
7n9TkLHHh2gVViZjAYTLJqpf+D0HAlxA9NAm1EWmk0SXLS3+1otKV5mr27nCan6sASLz0DRQQEs1
kNWcpFJ+doVQPD5TKXlF11PTZXyAMCPl4FHlCat8oX9G36Q4IldNSXPXjanbphuvWBcI3vNxHBmi
IHTRClHt9zJ465x7ZkTfezLQ9z5Rgg0g9xtcvelcD/Hure3il0Dobke4UI00Tnkk2tMKMq3+ettB
ooB3OrvtmbR6HXTk+tfWBrcI1WnPbuZoHvLUelagymGmgD6+L9G+NMTbwLVwHVUurysyxzhba+FF
ny2nb3qw4IlZEZQWP6HgQGyRw//E42sX11q8fjSfqIvnUsuUfbJDIq04NQBed/4Oiw8d1sNy6IcP
uiZR8IEAhA5MAJAvnpZQio0ZLALdDQs4Vffwj/tclAe3brhGc4Jt5gSvyScVA5eJriPYzxohJSAI
GxJaJeCN1i/iLT5U7YOiKdfHrPzmUE75HGOFewOZ91m15+k+g9/EtxuCLt59E9de+cTpar4GAZvr
dj1Typ0LxkRDHW5vIVbX7UTIg4qm44XyL76g+idi50H5hqjLKXhWo/iK2zbxerfqNskZkD0rIhqJ
SRLkxGuMVLQpQpR6V/sMuy50kk5fznvCamD4x8TPvHLY2m8z5x7p0SuYCujbXQgq4Xzyk0Ziqwl9
Iy87OzspAPcyDIpEGxIcAVVK79V7v9hkdHhD/HLanoUHjse8mnWzDhrJ2K0t47iMNuraTMHIwAKQ
dpVyNSvq/Os5TmK805HfpvjmoJVJe6eztHuxU0zE6tQUZ0J17vaduQZdHhA5MU2qfAreRJFOQQtw
VPl9HLGHW0qAxzgrgvrlXjGHVsQsx9o/6NWmj31sQpd0N/Zbpw1BJHrue6zMZ5Ya0qbPmFzqgmnY
603qFqu71hyLpjzQQL/v7//T/KLUm7BV7xJwyE/DLmbmOFu6Zprfdd/qZYb1cTxWfAA5cPskz4j6
hR5Q3BLu5W0fj22lpNZMiqYJJgFWpOwrJZf2bU9oF4XptNh4Rr3wmFTudRkax6qBpDWcegr/LKSv
B2lzrEc93mSd8KZegiJaR6aK3gi/zBj2uh0PH2zvZP/CewCHz6xtxX7Zj775R5kSYtekybCV0xnF
/xiHrRBOS8ha1sofbPIeebgnm19ekcrYAFbcLbtCw5Mo8AemY9SDiFvLZLftmWe4il/0dGtmODW7
wtTVanR8JpASkmKzhG4mtaBsuVyWspWuUKYsTxFLp3ryEd9Bn7oT8yYzdaS9W7sqqjwsf2HjaHN3
4wLagByIBBOFI9v9O/Us3LqFub/XTrHBxtDyWPe4bG3RfZoVDTfu47jf2sroOew6p7g+MN2ycN5w
jaAwkPEcS4bIzc8f79YwLtdXFxNcG3MAAmlxUjFdF6xm9/s/xMpXmUL5Ywoj1dKHGuCfrU54Ppnc
Us6jxIFOXzLgSEhublsNl3tYEhabEEZ8NYq3Ci3szkc+4LhNAJSyw6z7P16lo3vz3zQTlUPc4zrr
vRTFiaKSdDwMddu067niBB4pcgwg248KjO1aMwtEECTJnbnVAObZIvYfNuAzRnVCfSx/8XaT8wG+
y3L4Nt8qBkEhPWFDesS5caWIb+5730IO/WXXpmcXxCViARAQeZyUYv2l8wkY0CgmQqR+MDNDsT6y
o4Q3lCjjKWbUP6BaDB7cfpitfSL43xazXu2Nr3nssmAbZwz0lA+2QDyiysB/QeaDFsa7I/U9V6qY
RToJrUqXL0CU86hWjGBS9UfSQTkGCHiCcGNP4F8zyZUfflB0j4JJC3quMln1ouXFvsPJVNypmg9w
MGFhmVPqRidsU/5jG/DuaQmLogS7nzf1gjuy4EV6+HcQFQRHz/qtIwwfeT0a3DbxM1VABM2EWkFA
3s0+qGocs6FsHSvCmOgAMpSZfwN4tBEHgvgrRuA+CfTH8AlCXg8Y8jWB4n3egxmKW/WHdfpYnQgc
lK1m6FkEhEu2MR6lhGV1JEzOWxNe7lpp7zJBIw965oZRGSz6AnRpfTSAt2Msdkjm7x9S4zKkZmX7
uN8ZFpMhEl4ghP3ZPMt4T5u+PfNqflbs1qGt9uWuj2YN6bYkmzEt93n6snsrKWbN05VyNZF0zCG1
gk9UJ+39LQDFWA6NXhSNmrkYSeYi6MrsL9NKjacy83zvI1tvK9vfXDkNmtD0tHSz93Oa9jXZ5uun
0xJM3mipsBwC7q+Y2V3B1sRjqa+6YJdnVAijpJeFY4wssBaE392ZPCF0vRHQcf+a+YAFWu8F2KL2
ouV7wZyqbhsHOwlzR9nmphDcHCWRdUrj978YRNzNqdkWCfB38KcHOweR2SGs6hLHxtRIhDocMDkm
t5U226WtU0sGKTbV9iItOif3lUNlckZGX9TYkyM0vJsDsAiBcSG22UvbzmCB6O9Akmxv5OJ5vPgJ
eMO8ZlwmDJbWbpaHKWD7072l/bHC3E1K4Akjah4KNmCBue/PFSEP0Q0ZjytxtDp70Kv+wuFmGpdz
xAuf7Ew3kShWtumrrkTyZfT/WGGQLD7fpq8WOqroqAby8lMOiJfF0+RMUp51mELRcn4zhwXtvXMj
ETfaP2OrqrTDuJuCCpCo0cePOZwmqVT4ZIHmXULmD671rN8P3vAQBuOXUH6trtqmGFB2y0sFr2xQ
FkvRWD2iVOcIWZGeboDb7PA7Bwt9nHP/h6zC+6zYweBsU0zy2JQf5ya9ZZo1gHaEKLPSDGHjNsTF
CQXGvKlgfvrFuahpWyIhY5SqUzTCuH/hdo7b8B6+AmrcPE1BYxCCx6T9XLk7dq0WcijBdVMyyK4X
gcYPvpCU5VF8uqKtQrretagT6fA8RcJCZxUsXf7jw9FGT/JFBv4YllpctSCfVYatVUcigRG/aN6B
jeNAKQ7qotWl6UfbslaTeZcNnZYsDnh+zj5Su8dXsuIB4vnmFM/EolhQZv09jNvaG8UL/dyGkk1C
CdM3khNomVdCLRLyUEnyvH3H2HDMADfVMYQe2jetXEj8zC0YvDDOw0JsDJgeuFiz4v8e7a/OuGtX
384NxvyvA34Vu1K6aDWvmR13phEgrWVRzgdu6b1/iETUdgbi+ABMrV7HUtQgRx8R/RO8vIl2oLAo
obcK6YABkThzJLFDmWMuqjFCYijcIbfXLpm5P7Pn0RzOl3wgon7JqExPLSSet+oQ0i0JUev6vVHR
zheJ2g/5eOGIm6rKs9LXLNQPFU7m6J9KGxJEybApysVpRzeOlBLNJoySlX8jq95XhJx8h0Nw6Ifk
zU7fjqnSuh9Mva4oC/YM2UrozJpcUooFOFCyG+63T4s+K6mJjOWhcrh5VaBWlr5ymtLYiUwV+7rX
CxauC99QH1RzLZW5/7UiUIH1xPe9Wr1R+6ZK2fX3ZcyfBXWJbEi5Gu20AbP+GWPhsURZsTCv9/mB
pUcUUHlsv1NtzMD+d3nnIKdUJvDBhk5jZafAsikch5RVjRXE7zeYC1/EQpjgTfck2lYHPCa3CXSE
83l5VVn+jCnnG05+6U0S4WhX0jgBXNEoSX0BTNvF8zYQKeiu+hdAMw1H75L5lpcZu+VCfrmhwgnI
1DQYeIg8hVWIfxB1/JhdLzcWZDyqC8htGGacTOc0etDAAX59DpZzm168NLf0usobIX47It0VMav4
dUC4ZrDawPsaTWXT8a5Zb2tUbcG5BpJJguvPRkCGWzzFD74UgxVoXrxyG2KeHLhsm08zI7i7cp7H
Ae6TUDZde1xrv+ksVZuXWsILP+u76MyLbUBjfGWfQ/ZgYAu2d7tzNxtvNY49ZhYqrAE+iR2jkq1X
iO2bQx2yEHg2908XvfZDT5MyrAihumiU7JD0Uxs35GLsjzRz6ms+YSeiLprFPHiPF/8U2matZ7kS
cHtSquKYdDEHC1y/xczbQDN7amjUDeNf0blvAOj/uVgRhXH1bpTPA0j0k3yVnD0DJD/RQsLrKjYu
AXIK60DLx7TgVitLkW9TlQET+KzBJo+BtXehZUdg9M/7auMNV1gmLpNxIW0O7x7jdcAl/3fSM2L0
B0xtR2psStw1w/q5gOmHMNBLFr3CoX7oCGS53bVNSxw6CZ4FIofunxuMoFK+VyaFN2twd/gl7lR/
47hs3nwmbzXSmF7VyQpO65G1ox7quZjs8AnpVeRxzMRmB0AiIWlNnCepKPmECnQV89r+AwXMEXjh
rpXgF1eLEfz4RXKqrQr6Y3SZfm+PjDTHmqyLFqPhbRti2MbJ0y1wXuESZ+DnCCmCHzb+glzKRcaC
1uKV6y6UI5hA4HcBAj0ehrQ+iLBqazx1Xs3+evThMYZTj/VcT2yjaKtmEnhP2PCrkXwRMOSEzimI
AYNTiYaae0N8fFcv4F7QScvk9X1JyIQ/G3Xa+SspXqdtctX7H5KU0CipmyF3jcCSmnvDF4xG35W2
/wyW5YwOl37bZlCh/aYfdKTrDKI3k8WXAM/u3Y/uHx/9wXZtcSGnQCsiHHxVpXeafFwxbXfQMf9h
077YXaKz11ZLmLDuYEWPPt4ROxt0ohtiuHIasF4Ih36JL6AMFkqTtIAyxUhDCw3GfoD0Ac6RtzHJ
Xibj77NTmlP1FHF81HcmJxiICQu6TiJTVuxBDZ6M0TPHKufo7PKjbr0xnwD3Fry7d04Vc/GJ7hn8
3g9XBWGjkIf/oDVci2/xrXHaMax0z+ON5XsZEahU0aDuHbCIzSj+0XDvzSJ5RAtc8sV4xLoHbWcE
gZrTSGF0utFkGkxdJQ1akYvfOneCxP4Fo3OZeh6kuIn+eUq/eo973T8poPsWPLQujecdEQrkX46a
Yl8bc3i6GTLF6ppqR7+J9hmHvG+aH4lAN0QkYlr8HVn2Nu3mLo3iLrapn2ZV9Ov8zyW1ULApOg5w
zenLy4gm+xLtPAAk/qurufrfrnQohz/4h8G1UCYzBjt2GXMWLguL4S5eOob7WL68oQcdl31PFTKh
+HL2nXDlEd/JILsUY1wknPKUASeSIhJD/5KC03dz3JNib7ID6G3UcqWrva68C0LzwaPfz88m+e/T
mqOFCaAzwIn1GBKInQRjTQzyypjBI4wlCRyu5XFF9fhshqmeRNddnNaxpa1FvXvfenC7qxEP1PbW
7dzCmr12dmirySZVeFLvDZNd8kScQ5U4KFpdsniVxZlxEBpgQN75uzmrE36whakCicYiEtfzsb4W
qL9IOAfGcSEdEwXRiQPnUw4YExkaXydLNb7xr0ZcHV6PqPOK9imF1YZHlE5vTAMjqJC3PXT/+KFU
gNiJn9NdGym2WH31Mo6RpoPOAhpl5WWF+f4Ttet3FH6SoTX0J80JszR7OCqcr56DcaOEM+muGTHw
e3D7VkDHk69tdb9gmrnWmvs1cx32+QWBMXi+aesOpIvbVN9w/Ex5qXUym5OhmQDF5Lv9rq7Esn0G
tKAJFCKPXitU3wUXim2Y69C+T/MM7/IUA3ATdV5dE04k7RwK6mQEwanMW3aQ6aYizwY6y6s6VljY
lD1OtdDf5LppbuOTZsYsy1T+5Uv0VpLcQ4Ii4qFR+ndaCULMQelERe6joTvDnN+GIN1uL9ETTozQ
0qEYYAas949Yb+haD5VKH56eejnKRleoAwZObMCPeE9pjxaP358BgqpaUVKELzs1NEyJHaqFJR93
qD4rEgQjWDkgG3KVXFPxGAn2KFG5RcYn2kJ7lqTZ6M12SqxnWMAYGOnWvoh1ESOEmjg4TItVpXT2
DHwjSTjgskUIi/5/sxcwzJgD8N2tkysfJ4K0wRuAYacgTF/fnwgyEl56zuGmuIvQNrch1+6wcY/Y
leHuWw+DxHw+9ORQ1NEvQVac4/9KWHCGaAeW+c+JSmYalXY7tGLjZPHA90OLhL9BQ/QEuTdcfHPp
RVwl2ter+vq55j1Dr3RdjbMgkOiZkNt9IbIsGg86qm7YPa3V5Z9hjDIO26GqEZ8d1zQiEx7uCtwc
kaDqWB4RyJWIuYI310k6EzsYQ0nxUhfmBidpirXBntW4kM3GFY33KQ/Z3rXPzbRHdQMBkovl16PI
ntEf7Syg828FWwxx5XZVAotRTgUxIyW0nW6RFjfyizStoXkasOA+jYMffoyvNgpvLykYd5kWmyTz
55PgWE69ovTLKRLa//0LMoN+XYG9JvcaEt10VYounWdHj/YtCQomUeRVSx1DrvTwsvkqhUWb1vYT
h4ZFgtDOeVQwx4CDB/CtVkTIZ+PGM4ovR3CoifkGKqOJjzJYefXfK7FAL0JNvb/ErX8l2VAKlsFp
TQyJ0h7CaDh1kNxp97lkpGzovEVrdcxuBmGfm3oy7rBGGABeV6dGudoMkdi4Fo5LwwrIlk3f83mr
w0kULZeRz4WtyUnPb3659rnQK1flvx11f3QuFzkUZeX3hG15xz/2H9w62GU9u/gLXOZfJbflmiLK
2x9Bqaae+RyZYU3j+qA2NLpzLp8JIVjyZpNf9RNHf+K9O6Z3004jZ6RP4Sihs1Z+QwfOa5syGETi
ej/nHN6DTRZTMCpaBRVzW9bVlzZUOF4zncyzgGTIvpq/KtYzHBr287yhLTS4xGkdoE9nHq1LfUmb
3Y7toJw5AMpjddPiEN7dt9p5pQ7co9ag2aOvphFnS+cAnEN/Ay/fNSdpwP9nPyarGioQXnQIA49e
dC8mwX+G9OE1ov/aUvtKkzpmP3ZhzKLWujXOiU09jwctlWr5mPOwMczNm29PrVzXwfe1DbcYZlQX
TU4jzflpzcd9C5m5Y+J5jddeGDnwhEECHkgKeQtZQcAfQerBHJM78agyHys/1rSd8zoHYh834vbm
a60TZdcKuGIi3jrwVt7G2HZegxrxsVFEHnntNz98RtJFdZ6j7A1vvZoiuIDRwWdsvCi6nYCPIONK
DbgkyZhlAAdOeR9UjCV5mnSAya8ZI644a17fLcebwfWY86gDRYbzgkgltWr9/tTNfu3U//4ojZ/K
Mk62hlnyq3QxmdCFeiWNhDFVp9Mix3jkt+/T1/ZKKrLeOjhnLwE0xa4PYhUZTcSrXDTNbxROe5l5
hJyXdHuyqWLcNU6V8VtTpKmar/BvWI4m6Kjxlipx0MpNl179i1m6MQkncGWSQJgKmqyv5c9c18N/
PWTtEGfANpo6rF0cwAX5M27r0YSCyaCJISuyt8P8M4ldSJK503pU0EMl3t0oE4Rz9B23GaSK23bD
lLCnex7M5JUgXeDQVPm1j0q93kLmMgmotMw8q2RPE1DaIVWXY/VTUlWpi5ZqSz81tTqK1WTxigIg
6D1FafycdbI2gGbL6oU3QlVCr9TNyEj6Ve49Ux61Yzn7g9I4JUS5wCmi6rpu5lfwgCN1ijhMJ6KP
aPf9cYxIBz3oWQ9dvqjRcvRhKfxGOLN1ERsb2QN9ZWl1aGY7sPDhLrhq0heGJtkxmtdFF0rtI7ek
olfEselovhI8zfY4n2Dhen4Vm8ITRWSPFnRw1Cai7uW0zbmmN65v0CzJ/hiQZXyowoiI5FEzLtB+
i71iQJf603mf+kiYoIeQAFinZQYiqHyaDDTBQWrKDiCQsP4aa8OewHpXoKQi1eb1JTKlvv9apJHM
hZxpdRZavI0h1qlt/HYeaF/nr7cVWw2xccAPR4HVY4DdtlMxoQY3bg4/hGy01behhNscTL0FsnVA
Hh/P0JjwyMI+pUsewgL0Jv8xvDtXV83+7HPXBJBCo7EA8MRfyAOc1Fuf93s/4POUK8Ii6pPuOZ70
PBoAR6RvtxYf2OXwE6o7XqxY9DaoGGWbNGDH0t+y/Rny4nelt6vjYPebYzz5SLxwSTlZPAbqYd/U
aHCuVefc6TKJ24l3gFcnayjAUxw/fgIxh+BIReEwMjvboQTSJKZ9/9UMEWye+yAxuL5clIimYyvW
xNlgw+epxr4xgUJZy7P+795IixY1ixUzrWZvA+E3q6RbM7oFy+5sqlzFKS7FUH7jph14B7oBvJtJ
lkosEEu0/hfAJJXVTHuRRFQQKGDYJzqIerLUIno162p8aKznin50KEGgUbSdLVz++feTi2Wie7Lw
SCNVZEHAoIbwp0BQ2q9cEqwjZEbtBXQCkQNpkgrhGmcUT0Gj/4PTi5wiPYnn3a9YCdihXduBlbiY
sYvz8kcH5ILfuUWXH/aWDdzjIGN6/j4xJ9FSnSkB+nyVt0ULc3DO8gRMtlw+jSCU/B31+StAozBr
E+6iaUCW2Z5LyhKaQzQjNUxjcL+geN0f7PSSvBLUzQTLiQB48OQaaIFVOBl0dIwnrB+eiNIWSDiA
KaTN4asV7acJhd/f6CHOEwYDCVnMHjANw9NqfM3Ps8EF+7WAnmY3YPzcSULgv2Sv6EZSThlHVxxc
DN8OTC543M64YiA7cOVLuM1b9N21cm9MSMrV9xrPnrA6alAWvspnvT2AHQDPhNgbhgPwESw9NUUb
ViKI52WINSIgqTLsUkVbKE+0z/2AlRZSVghk6bgDHQDKEwfWp3JbJNG3gcUidfzvHuKypuD+3foE
tnRYZo71vrFhHFDSZW5Ajn8hrbtfRwGc3eDbJxsSLtY1dk3sEOPQNmdQGO/OY1Ej2YeG3ULZo8cA
V4XAdhDVKB70W7edX0bx8UrG98Ri94HJS/VYrnkH7GbwHy7gE4kVmBR7vixlU76UyApWr5I3+JMz
Y4hqNZNTjxa+vLEblARYuV+m/0CKTMi9eQmQED/JdSVeml8fpD/g4/e/fJruxtE1MLGaxNyDasC6
M+AuaeLpAQteMQGOTC8EXSu8lC6fPE7r1EVoKRo6qTHt4c1hzA3scTXhQU2nFb0dBvV+O4lYPSAc
7TMWRmxm7Y5VVXKGwAMEt+mxDCo3h7wvaJ4s06mKtwtJQ5pqXWY7b+LpqtPruv4yEwswIBxaWIWy
IvT8ll9rWDdRHbnhcNjB4Ag8/wsvdKKjRZNiHYZrrNyEtwD9wf81leeztWSbqInf5Cp+PLVlste9
Huh0mn37r6MDaB0Slf7ZVpceNTPur/KsNpBMFf/pIuVAPm7m2bn7/ghR9yQVYmpeuqCGHAN6pgL1
cBIpZHCZpdz4gUbV8AoEhKD1zJKvy9Z1xrONKF3oAcVf4aA8n5KYcvMzHTFOodZ42J+84URTFh9q
a2+9usJlv970t41QRhfKFwrBLUWgquBcFbmjcZJt/aPYOFVCclEaYl3349HOzwVQERUZNE+55I7g
P9I9u+k/JX+IXtSWlc6Ad7qkSi1dTkS5zjrhgbB02MkcQ5ay/G4YiRuR26e7YnnRBhN6sm7y9k3/
YCMRUOX+K3pzU3YCayAV9fNtcqnx6XW4aALNQew5CLrFVIpQvkpJTn31TJ//0VbG/ZMZ2tjlF8R7
35aR9YqlNsEt99OfonIFBzB4JlfFDwR/ONt+6CiyNfDUQt8fnf5ZoEhODbC/CgISEtAL9uvHtRRG
7QSFBxmLXovfA4W3JzKZ4YdjPpXjxt9YyyQOaX8q+y3crD+eE1WXc2xqZtiqdJ0b1+Yja2JEj72x
00q4dWJovxCFZkT7YyJpxbjGav9ps7FBUVwHsl6LvkLxJKQpkqf/GeOGc/ynVZUanuW75MLFWQ7L
jINlHOXoMCJ1UqlgD6T95ilnrL9l1VArExD+KQJXj1TiBGUVTq0Ib59fmeOAHMhbZ3wMM8ncYLV1
cf/e8MsWtOM0wvQ0wQ/xy8j5RtmddS08iaxUen+lJc3nBxsAkE97PzAyIXoh3s0NpOA78OnembwQ
cT3WuREi6CBsdo6PE11IV32AAJsH8cPPGsgQcFo4ZPLCC8lJwaax7kkt43de4fiM9tO5Qepo0ASd
AtbcqMAj6cNBBEvTQNNaaIRFHraVY5MQVnFstckhf3UynHMOwvkpDFUKb6U3DeDtbHr0TrWmQx5p
2viLz7VppzKD+vCmxPshQJfWrfO0RQTOfDKFkOu88bLACtpZYeE3422Wmc1iT7YA2mimTASHKJjV
7gUqXlSivJDFr3ZSEra6wfQrKE23H2KEndy4V93qteDr+s61oRk789wcyrZMVY2VfZiJEBmoko7p
07I09SjamFCoWr/fuNxeugFujFm3YA6spYpy9yLdVxGoX/TVgOpbBWO3KYz91NQJThJb7nPB6YMx
lHh0gL5o0VfDfoPGRh2YA1KRl7QKhn2Yqmp5sMd9zwZL5wP3RrCTC6gAAKmUJfLwtf09udd5qjht
NdiMxFUQ17JZaXoqJdDEnMM9Lr4+BZDT4ezQvspK8+vSXw4XAlpZS0a8gLjGrUh3sjg3hClregwO
jpciDnS/b15EhkU76AToyK3S2+cwydNAISL2p39wCk2Y+5f+BC96ajAX+eiM8uqA6qpVeWUgN4Nz
LttO9Kb4vJEL9CaWYONlAuzOpdOAZ4tJd7UtVA21Jo+N61i6jlnNKMmxNJ6bc0XgASdMsi6HilR5
PiMbuFCq2HwLG5TJBclEfFl/zhagJ/PDo2SvfEfgbaq0HQOqXo62eTF2Bt3XjmMk4y50hFup/q7b
8R/ISRPMpuSzxW/+BgITf1TnxCzDT5Nc231DcAk9bVzjiyEQc6Xk3t+JuHvzfm0QRYHzB/X7N3IN
/ar29LoOIKwEoV/3+tjUBq0R8RIBvbGHy5cSO0EYeRFCYqkRqn8YNkeDP018TsKTls8gEcim28JY
rTrqeNNPUSg9I7SUcHm5S+PMIvc/ygePzC9BZ4AARSaDYC6HftOsOai9X0gINg+CQwurQUBsZway
uTcnjCJKTpnen6qMlVek7PSyH6tRoB3Ufq1fXE9ughifp+QfcWDRMbqBHgszIK5DBAFi6DR3ElQm
ipOUIz0+PTVAQBk5uEkWKDgJrOzsWfj4C2p1iWp9Gl+jJkFVNh1ykUW+qI+hhXRFFhFJly3Q6wuI
CSYq5t/LFPEiE2UnegyCBtQavdJjRt/y41C2oc9V7eiTUfPV018+9XbfWSMkncXr1LvRxF00lTjY
RQ996OAS3kDYvvy1/BXZMvUv16HU8JXtQwvFRaOqR3y91Vhdey6igaAG0+JQs5ojU8vDeXnSqfP5
QONiNJ4xePQBogoorMwnv+4r8mpsW+iEZS/OR+OCfo1wE1/9wZqrF0Bf74up1B+zZhsy3z2PwwsL
JPRR9QehmF2loyaIptKfYFiCVOdqjnO6H6mwywMGxoNtqvH8masWtZDk84oeCxw+QRrgn9bAHsgN
xu/1Lx9Q6Lr0Fyn8XyTwSQa9kRZ0A/GtdrS5VPlk0z3oBjQwVt3pygCMGIiRv5gXqVLfu0bn7aR1
frY6kCKpd4PDo4zjXQaCgP4/KLgwZgfMnVQFUoY0FgX77cqrb1Gy/hT9z19HagsCWgbTywTXT84v
YbTxFXZW7RnZH6v1V60LKxwsnC3ajnsBPcTHH2lOkPzgQ09VjKcYXqz6piRx84AIkTc2fQrXIPjz
DjHzGaBGqXBIYC6wLexoRBu/yfTqrqT7tIKFx/ooJnUPWGaN3TORP4aLf7bCoX+REi5T1MBM5M/R
yPqDKXOoBpd2MiVc3tG5q69YwfMIy6SySidpiIWlEv0z4DVuXo/pLuTopdDQXuxHLbXmr+lNlIx/
++KUwr+68VIfmFkhKVRTfY2Pr7YL/xnhe4h/fqIEWB/POdPPDIUIY5ofGdMchdfAVNef4ynTDjUa
bb+kyiZmQSdmFDZ8KXBV1Ry++zwJ3BMpFCP+q/MyP1vNgdnaukgnEC6p/mtyVGg+1FEipv/e6Jwc
uZPeaAgM1dLXJVl1HXOILLgY6C7SyiJq3uPHBOk0f5FPZWVlqZbDQHGA1EXQmH0XZmgNqjHQOv1c
P8E5yqMQ9kU2yUipNKyBRaM4ZzMXGIBFzNTAe8gFbnQo4ZuBhFfdul6yHZynzKIUfNFYDyVy0s0h
5zH2+Rq+KXtZze/DMTNi3axddu1QguWx9SNzZbDHDyTWZ6nJJVUIyoPI3svQT+FS+qOFXJb8UgOP
15xDKsTQKW5Ig29hSaq49Y91HJJLQz7k0zoG0K8m2gfW0QbtEvfrZuMD/r2LkNNkqElZYboZ6x8O
thM8h9Y1qppGoJeItl6PDgfuZh1xR6Q7fEnemfRAarhaVO0RBi2SKEImdXFgWtgyL5LiIva3LHFC
DnM430ncBIV6+sGLcO4ec4Xz17cohEyF7Jyfxev7x+VwFeJtfpSme8O/+EDMnYxvwqyA+H5TSz0e
ulIsZW7qSOtq1nK33W6SsZiUYihk9E9jVZJFGnjdnAe0v2abpMulzzo8NWgmwEg49g6ncuuuRf5R
/T7iIGSxJ0/2UfZVPjhqiBgWx3l0uzEPFJQXFl+0X4KAbEVjZEMEXO/iOwKr6/Nn8rWWfTLpeUca
PMecdHmhemxqNwXRq+jsZhWiJK9OrDojYExePQyafhD1PhJKcghT00y9jBuxnaztOH0qXZ+PIA/i
85YWCCwphs0Lci3jZKrvqmsCEwDrWWsLv1NxAxcPD3TmZSz6HoyN0HDSVvJnlQRvS5B0CnaHaHU8
eyRytepFW8o7z1Jkx/BLFPboxpG2ABiQiuxtYENHdnHIRkYXcsJXVL1CWiQyB/ggTXXA51HNLSRx
h7zdhRl+/J3KT3w0+QAP5TEUVdP1DSTmemaK4nrobGRr6C7j5X/y3Qv1nyRnYxaPsdMrlRE7Nylm
7QjC8fDPqc+erozmQqz47ohcU2+rRZKAhFT1OBuKOWIiixc4PUkzWm+bjy0eODs1ZLyST5ZQpbkw
azwEGyHBCRS6dvnXtfcwxW8/bBQJhDQsEmEozzNxt+Fg5BY7nIXbl38BWppWVmpfAai4VPPcMn5R
/+Q5xYdTRngOreT3NBae5CV47Vv4qVkkpSzwwk+AT+30wcKz99ER6cGmLrrsYklmcnWQmUdHxV6/
Sc4IiTUlIJT4zmf03u7kwy5Ki1fmMX5TrRx0NaI6gUiN/yP7UtNXonEDlBAd6mRT2AcP6J+FoIb5
fu48MfA8M2DTw4tQtbQV2UIXHbMdFtxrlGC15rejomzFwp4JthyYam5nYWbPfNIxEOJNCrP9wlad
WDkJs8lor1JGav0SizQUYWL4FVjugFvSdi2zwNFlN/aKqToCLW0wurEZt6WK8q6zAFZyAt60GofQ
d3nuVuxM0Eg0p9P/D24fo8ymMofEWWiA/5MZDCTeeJFkGsRlbPRWRIgq6Mhrn2+2c84tuc7KHViC
OlzLVRFCoCL6sUpAjLKNJCOESHxcsw4V7I7cDBtze4qNGP+I8FeH0a2RnhORUL+894PVa8ClzOiU
4OzYAED6P1wEmC8M6BVh9ztiBE6IqTOAxaoSFeewy+Q8K9ELKH8itwXYcrEC1U9rvkV8GJS+cSQH
Tjh9sOCB6KH7TgJYqoEkgJ1VCuopiPRQRwKwTm5QWjFLE8Enzg+LGRGP6rOXLGaZH0mnTZ2ZRWG2
ynS5gdrCj3gbFlFZFuosXVNO1waIaJO67v9D/1xXPq0C7scGWGc7NZSb2pxAidUg8/ZIryl6qWV/
AZIQz3O5XxLGqdEiQN0AyktrRxY6H73OrTCaK7YJbyRzK5lFewjWw+DCdJRzn3DAl8mlMGvfLJHv
nLZZIRWxhanMTVmhTEW2mWHR6EzzYKYHm6/6AbmMrSgIeryRyZhME4j4G9dAuVXIh8t/G0Eg4Kgp
MbDBajzf0bL7s8p2TTF+9ALCdsadHfBafcmTLm+Ce33Y0Zb5ja1mSUUrb4IvdZYWgpIoLJeV7t32
+/KJMSHsXTvF2Cn60weyLgaRy5RxPaKvW1OLzLRSp87y9ZHbPeR5ch3qLjxt5MVjEdv/M4vg4teU
0u6kjoYjy6K5GPiE0Xcd1iJv1Re7UKs7P0BH04KWicNiHLW8JwO5cKZHTZqhOIxd4sYVXwSMUMiy
PB/npNXji91Dsvu5u/bzEZBWYKSoAl35o0iV57vLO8YoisfUZ/dkIBAg+HHLfp9Uy0uwQ74yJejo
j0d8uXl022cq6daQxjZ3nsTbqKBzeJ8BMgP9hE8OEGzKjUp1pC3ealmy4rTYyRL50Wvox99cxvz6
VNOcMDiemHmvTfYgz6SXW6aeir5jN0WAkmyWJfyjXGv8NvzT9xEmx6OEiCqjF6UnvcpmaLzanVDu
Wxch9HiGQ/1dtta/bl74HO+BISFdtDqdNAZMthzDC7w6JZrnXGJFPf6zU8GNuuJcGxQNGXaq4t1l
Bun3FBvzHPeOQD3AmrBtH+/fkpHZZ/eFxVIn5IyYCEP4aiZyN1k9vSX4z2NGGyA+ZTH5s//vDQWx
D1PmhPPS2rnDcO8sXSNNFFRnb10JoChEMISg1/EK1R4WPGgvh39wwcKXLFRt/dP9C6G/DwQKfcWK
cBoN8aSsu8jy728k36JcgRGHrREqOhQhd3q5ar/xnROMkZAH4jQ/umCeY/dM+BqYMZsqV3der725
39ErBH6cysvoLgI0YjRiVG6yESzOKYR/5mEbooDIe03Cg9vWRZifualCJp1ukcpOs/FztOPBdgsh
KHDtFqZGFMYM2Mi/dZM0C85sYBKJuP+mz8KaOyTx4GpnP++DUq0BCG56vS6zMEu9iVOui6O5edLK
Il2eE6lBATars50T/CupdQHkiuJu1BYSr0KO+dyDsxhshh3oeqNlXxaWcM7TJxJ0wx55JZnGne/4
YTiQRA3bMLQEQTJZituzC3rEuK30ofu5mz5n81qH/dkdsvgpZwH7VuDyor6fKTs8qcogQFpK308F
PX4G4pxjJ7BAhi9jSONerglg1iu7TM8Zov1e9ddbNDRcsM2SEf7oqmeXl9TkVG8icBGLXwIqi1/5
xFPDrEICCj58NgWoT6xABs93GjpgMiR3tPBKsJE2Wk20rcGH63TrJWA0UkimZoZx5nMTaogiRiHk
+UQiuf8pi1RUTxZ4Xq5p+hi/egFV5RoRp0C8X3AaoYp7gKkqv524OCSZmIu2q58SlZbysHlaYrQL
1eVv1WhBrUTwMi4OSWD+fCWLHac0/JFZpjT5F0RUpzNYb9bJCyg7IPuzElfPfjJ3l5Zu4DKsDFAi
tp6COzNTUhkuIV+hl067mk4Q/2kAasZVRIqOxbrsYi88f/DoxFadOXmQNdUYTFLpYvzeVoI85n1f
9yZ2gInibxsSKEEQMgj2a3yx5NRWkmSvocJfk9ce5zKgcVzDC8KePQNrR3wWAUhmO40/rbmRHzZs
V3OmiWVtY6/6SJXfbBLc6sbto096RYNECDShkBK0MRdW0c/NugpXByeaE2EUH1M0SZdl1hcEhGtU
G1m7Mx4Ok5JJFcIT6GTHI11RhknJVGRylH8JmqLxQaYr+gQeBJVzbMOwlC0q1nTmgfeRK3RbfH81
NiYvUFtHzU47t80DArbvnaRw2ofKflziauRG69YZ6qf3N2bH/EcfjJpbp6yy6FToWphfRp7sFOFo
Py8ADkOJxp6cVk/mfHGT3eNFpN6dJ2AzsBMmZWobgUc640cjHu47ocjpTFVYR7IFDAZz223V6XAJ
rH0+zsy+yOL5M6zzVxZlkBx4zbAPeFKj23tKdGmBqlBLfazjGwVQF3POMGCnIhEqZp2abzUJefdm
TTohRcJ2vz05hX8jkXxCKZq1uJz/P/B73sGetxlWcr5d4/bNm04b0Mjy2uYKgRT+rhBIbDDp0K0v
XP5upd+JuJIw9LEC3JNLf8d/vVHZwMXez9JUwoNme2sNzOa0H8xo7mGuV2h26xnDyn04ZZwRZ13r
5T/vpCvd7iBBca0NM5aSIfUcghMDb8QQm/UuCDiK62SIq5IS8ziXhhUJTEcVul9KwsOf17CTrf9C
jNt1SFkx7ET/hr/s0lHLbuD1PMqPgwQvvZfzc0mjOLmb9ndSAgi9c6GUe6Lr3T8nhIchdxC0F9iI
dqqciLW8blIA+ZLidu8IqZMaz2lUQCOqF8rWNtfq675cHAb8/K4r5vRvbfW5y4YARtcZawdyScKj
t9m3H9K/02UINp/P8bFlR3k/G/yvlRQ5PHSHQExFcCu+090ntmoByN6t2Svg+Ey/z3onC+mqWg2P
lUorAPnld4Y0jwWQrwZvLijvVL7et6BZKzKwI9EEjiAZXpnkTm8GsyZbBOXVINTQInK4j9jgp8KM
g6eyEkMql4R72yi26OqQoJhjkXYekUQmBZEAxmK2NPF2QZVGmmv3HUEH7NLyb7w/Lx8GOBKDyJcg
8SIVVh7gJzOy5oH19M9SxLaPLBeTUpGdIqiL4n4C7wVF7Svt/9MW/VLe5iNEPesJlFi5NnUTihT4
yR+IqpbNyiPrphJPzfrh8jI02bNESOMgIbQBkDbx/IzAUDGf0X8Cd18AN2O4TaTqNAtvEjgvypL0
Wz1/Vzv50VIliaprCUadw7h75f7F9AM8PsiQztItUBO58Phm3gmgWXzDP0ghR6iNnLjvbtELpLqd
UICCp8Hp4siNUcCKkqwwFk26hmDmlYOBpLwaiSBUlWJ4tcc2w8+1BTHyTUn8GcQyGM6Wisbnhd1H
gMyPkUoQRgEh+VXMzJFasAPq26++mW7RvlUYOeEfkehKdDTHDFIX2x/hhFChRSOb4YlTZnTegJku
fmOz7wY99C2SwCtXeYZ+gKw6RoICfFhmlvEM9SCe55uh1cyWY+MqJ8EeBX0Puq4r0bdwxOViSJDY
4H5RddeIsvTAfyIXnrgf8rf17ePjdsDVy1RAeyM5htuxp7wZ3EXGd3ilV8+Kd9g8NNmFhJzjL4Yx
D6nw/8pf0qRHqYbbpqIE3ETE3QBFmSUDbUbqaR9Obtq85/4nS9yGB6TBJBdjKN2iQ2UZFDVYyS8c
b7P3yCSsqzOcsGFDqsAucyzv2gpJ4dvCGbmKB6cOpPYkS3kv58gvpL7EvJohO7x25gcoamJUKVW9
fHc2cHea2+1vZBGQvPy4ESA1z21lAwz0HhHawfJ1PiuLlPzfFPbp8dZjKqI9a9/5PdO7JVNQnpb0
61fwZo3sqGzKZm17LvtLf9Q8GSM/d7aFOPvS7/USm153hOA22GcfRghBY+KtoTP/gD0/qGoYLEd3
ADkbkpaPfXl4k34YjLbX6Q/b6sTsyThzBricPqxKErIRWDrSxaYZBl+hkjPySMi0L8a+tfzf3UDl
tz8AlkcB0BbKDp/zo2Du8fT3TCQorCMwsUNk7iBWRtnCZOTMnBOmF1LO47VBBeNR/rq8sqgvHBrz
fPYEWTiV75Odejy1NoNKwrY7a7tSygRnP2fLnYDZty2Y11Ap84+8Sbx0RL8rVb4olR4cHvuGvOxK
TWbnoAe0j4LYdphrV23edK820rJkiY9wg+FjmPVrqNmGbtkiiIEeG2pav1k9GPeI0XFQJr4fslg3
SXy9U20PM9yo06kNEv/ABczCyyA8THAq2GNtU9Xu43/HxWPQjzlo+kPHPeFy01Bd57ODo2VKaJ6m
gf9MhxnipaUA5AEGDgAmKFZu+LNEeMWtVeEFFeeJoNMGkRiZ/w3YPZYVPIS3+1gH8GDqu+y/EPJw
248ax4cTwiL/q9DGLi6kcJCfJ8LUuGFBztH1cR1MdHBb+10VfcJ4EXyjEQqGIdApXHcR4P4TR2B/
1aQxYUestmch76+BkjkHGl9W7yjgm3I6ef7DNZIXSNly3AkX0DbNyDJKhnvWXDC0D2kXl9QKtJcm
YYz2dtOVWCthuH6QW3nrl12isfgT7+ht4izPAr2TVpovbopm2ApQH6kQEYH7DrOyAQO3eatfporW
kApnNpfLfRDK+IIhHNVzj65lCTZzrjw0UxymBYomHir9O8356faU+ObKzl70wPcTyS3mWj6IY5MZ
ZJLwJXxa0yrdwgOnsKPr4YldcixR77tmPn1Wtj0Wd5h+RFn230nCocBDTxL3NcySZ90mS0x5O5Kn
T0OU6lRES+fujXt+pk4XBYjOj77zUsXsVG0KKk9jhuLMh69IvEAcP3yJa9P2aOJ2B0lqeZ6zIi5E
fyVVEtX7JXFuyxJv06IwdUd4/RJ14J34KoLa2n3h588K+FU+qCtMcSOgwEq9TqCtmx4RaL/U/2Rl
4LjR4smSV1MpLLEgTKkXDpThQcuimQpFHMN0Dk7C0XJ1qy3HqSpJqYuOx9P0c10LQ3Oz/B4rr/Wa
2kgjh53rwHkc+nb992NjY1kmoomM+/sPhutHJJNk/dfe09J026nQoAT0d4r2iG/jQRy7wdp6ZJ4g
4xS6pb1cTqcUxJTefwP759lvygASbaCKBBBqE3ClCj+blc7en2N2UBC1HoRV1Y8pR2lEsDeTbyWI
nWKmC1LrDoHJlQLX3tlDc+CSQ4luMDxigragfqymsxDH4oQdQbhcOmCoYHsesPaY0qEneR0zvt+8
470d6JNuMqEt3IShavvL8EHaMGkTEK6G6vYkMoBowS1qC6WdVgQ3snGV/xUrpQXxXzslhCQ6gjUW
eBRHwNpdwsMICCfL/SeqFpYRIy7n4/PBCvvHCp1iAJos7ivGzch1ur8e8JQDL2sUOX7SRwc5AAY/
yX2r5CdrZ+KU34L65XgwP0xMkpjF8au6RQ6I8YD5NHj106V54LyFaYb19tNIkGEVTP7T1umtiEzZ
kcSC3hfJhYRbmKs5t3Uaft3yFXyVNr852iUY0eVAajBwghvS4aVkrJI1ZVrWoHaNjtLuGE1/Xict
FjUlRYiFCn7fy1EFQXxDlDnd2UBv/R//+FvTD2MirGI12UYCT4y5aOnXVauVZz949O2UPbzpl9Zp
qq4v/HNsO7FuCOr2cLpCQzKkFFefGCy+4pu8vMi/lza/ExI4R5mwhce3+9pGq1Xzqb/cIN3ruRLw
qjbZj9wl0HkfOAKONSuM/Sj6nrgZHFx5G6O4U5wHREGLyaQPJXE9xZdRsX/JXYCiFR4inm6iAqkE
7YS9njoYk+Z7aDnZ4rj4jKl5H82KTQs3V3UxP7t6M5TQrHLvOdrkF1blIrNKXdeUV6tryY2yBcUL
kETTnyGnI3IZQ405rA+BmT9qApuehcJB3VUgU8VQ06zdLn01BGoMejaJptr8vHcd/yESm80SMdbK
vZQ/L904lsuDX+t989XwsSeGdJzyVxVQGDRle0QUdgaYgdEejBgnDzHhcJ9RdDpNHcnv7z215IzI
/n2R1B5SE67oFrGSNVI4DXn0HkyQ9KkXNvzAjzxtYjDtD+Kd5pZoB0rowvJl32i3Klg/3FFdChhG
mqbv6inTOm2UnACPHumdNlADZu9yOcuszvxpJLvx4sm0UdQsXrFA4CJQp/RpGG7OYtBqFDeZlJdz
FXKf+DTbVePt5u4zs4+ZCZxgt7+rJVLII01lSnb8/IthPaLTMn4kBJkEHd3KfBziwzS/s/ix+P8l
ZeL5XkSOuHXRpIkaA0Od3cZanCVCToAq3ppGBKPurVljdbQlv4dg9ck5RS3uNOceG8VoBYm/7HbB
Nx1HYKC8JX1pO6JDX9tyt2xLOAYywaUl9c4VslVZ4X/6scESbVUcIUzr5sKUtyX/XQrJjbE8WRM4
ThW4aOkctkFOX9yqA9Guqx3Qm7KA4RMuDnLPyEGKh+YndpR9786/SmHiVAQZyQS70M/jFRkrxlfv
jK05WvYkMH+2Oz5iepV2jzuq/1srBChSTtAFYDCMoUbzU7NS/Rexnw2DfelUy7gbIow+em3byxQ1
iT4nYW19rkiOWAHbA+a0LdU+5/FwRTd6Buob+vwrX2u4/sptovK7/57uyWCJUYRmnI1THBZ2PW7L
iR8AZlij7Ab7YkM3dYhuznnqCo44KowdcD9FhHrMtaZypr7FgT/iCbARDaBx1t/oiIVgM1LFB/v7
0dddpPT3AUbLrNf4vXROTmEz7s++akCzkL5a0wGMfil4FUqqtL6bSAZ4OLzJsH3kkoOWmApyng4P
QBhtukRTRNUc2Th+V+/wFepQS61TXosmo/V77yDQX4afSH11BTqWK3yI5goJlBvuOLj14FurUba3
pRoaHTe4gP7lIFyHRDkp9OCRx2wBFIR4URXi7fSXay8FA8bU6ga8IyzRqRFSnz7MoBB1EecVwOQQ
1bgGR65gVvPMPrxpYiX7Dg1BHY3TS0Sr8DbiV5j3TrO728g7qvCvpqMTopu9fkBb3NKGA+3h6zGw
pTQU1nRPbM3sfbcVeeiGA67UgqzCqHRij68w8gmxT2nqmDS+T0eP25qwoCinn6nwpqZGlviiGAci
t+E3hJzDz+LYJYokQvFX5zsPl3+rJkMLGRa2k2qq8uYnYvQV7S+T6afCiqFf5nyARIxhVF294Vk8
m1DDCXkANCBuYGdn2tbXAIgiThmQyVZtdqbJRUqMxb65E3zGtDcy5knEeysOSs0qmMI+IQxh9NI/
+Xjh67LQgMOhIVPQVKOpEotGwTaFg54hs/G+XcMdpHAmdxvCH9M3CO3UKwhMlgcUyApPpZpdS8IY
gltPVfkxxTUGeTuO1cOgDOUKkRXP+iY5cfK6bqynD7WqHFWXQQFODG5FgvEdU2WET5SinkXQM4QG
rMsbuJ0HJBibf1+ElVr/I7O1glCDAz9/NM0xxsJlSYaqLosi18DskqhnopasEOYYbG9bS2Pg6ce3
xfP9V5uEn3lnMh6FN8Tl6bRlkJ3w/5xJAsM8KYQGagNzHzudaySH6AnzwcVbqMfW69edIJKlsS4L
wgV036K58A9KjhFawukgXnWoybYs7dxm3QUHMmrg5JZkdxldPyZYzE8jh9GQcgCKb/J4nlyuf/nz
5+2QtTzMqa+No2ALlB+tEBM7Fq/qjB0RTEspNdvfg7DI6m6OaJLdCirkDm2crOnvlfnyV9cH3o8u
FZyFJtvg9BHOyHlsbvSzPtqXrPdwlYFRn2iUYxGH/RDp6u8yHkVcGH5kiH13sglFnLGLRG8jbMDx
Ya2dYhZs5i9xzC8cxWeiRAKwYhTweIzpA+bn3c7MF7WpyQh/OwYdgLLkM6shfrDJscAxGUPMTKbu
25L8qZP31buYuFwLw3DXYKZDbPx6OvyYDg26Qy5ZvNpvwGoVW3GUOxmKSlZekiRcc7ZmDHWpOhcW
k5X4gpH+vAdqKJmI3OEaQSvY6jXV73zdG5GDNGGj7AIx0RLx3pFW+sXFMjBRW0rco+wND73bDjQI
xjyxfMOMb3/fw4UxsYG0VPGhYohrZMB00Z8j7nh5cusUEb3fFUy4LceLQzuiN8pxSYcddGrzcWxI
r8PcPlM0CcfszsVzq7Pe7wNJCfWUQld7GjMLJj+ldSGPXyihNBT7TK/VvOOh0C0KcNXk1A7VAslm
P6hZzE9ome5jXugLnbtBbyEMW9E6QzT7pAfyyllNrIkk/nr+Nqls4GaQbEJZG+XVAXaNUNaOOY3Y
neZyey/rNoqOq9sCayyZ/ASHmJzITw31eY6tuOY+K+c8lic594sjmCHcCoidWS4BNel0Nd2ognlC
ZrPDHuxRddkfcootxL1rgGGQ5k2YOg/Mmse8/WceKwZ5/oqI5yY1aoodb06iFoXmSVj4trQYMewQ
fyMjAg4VBhcHqfwAFQB4ZiGLeA0F858JnQvAG5KwFZK8UWua+nPyuSqcuZp/8/0/apyDb5uOmopW
xWzBIGNwkL4d+m6Q7bQvaIA2OIFz87fX+vh3mjpWGdK3G5xfI5b22yrp91hrQM/gYew0Gd7RD1K2
xe5/JWikdkC7nnr2BCxiJZq4dhSwtWYLENrwRhbUAAUg2hptJMezFQE5MFITEfTa3YLfWezKpuFM
cFyFiIimtfuxh9LlX8/fz4ExQm7pqti0svOnToNblqmdxF5/sueY1eTfYaKU2s1hLTKgWsH3qc+2
CqEBhFRS/rG5Uvwo6n2ySzLF0EFMgHC3YibKYzkAXOyaKdb2O1Yt38pu5TnrtfatuPFv+oj3Dx/+
DkR1XNGYi5s/fiX/nDql0wobcm5CMY6oyYk03Dd3GGDzk8f0qLk43HngTzeYZdtpKI6xCU0r31Dl
twPmwIbQ5B8CZTjJiYghtPB/G0acJul696nvcqBIqRX0bYjcoG3PW7AbAOlv1u5La3toq8QbzBmk
rAZqMye7M0VAWBL7Uo2mO6TZxLGeID8x6rN++gpypeDQBZUgpbGWs2fuFYw6fzy/lk/Nz1g1Clk0
FLja2qvnbOfi7vXii15f+szUyhHk5fdqQEfWf6is7Ig6TGxnDVJ6AH/IUomEPJnEwzLTrx0sfN8o
C9J9Ub4JQBAYPG5od3LekXMsISGLVntu9eZUzWN1cZm63mVplIndmonQB2nKYLQ/emzeHqFIWCiR
LAadL853FJnuxcBfb2EBsmFS7T1WzgD31qymYJArro4SpdTfRhi09E4CtIuSUxU2+V5BI5pSJYv7
qlJCJlzst1EfCvKLyXeaEr9fv1reM3dYgt0aynd7PhKFWYG0ak2mn0LboE2MnLSXj1hkmjOVra4+
VLDZMU8jvwn58Iwg3PeYereDdR178l9fMzPKqgHQqpu8u8a9RBqkVXoxFH0wecBvgOxkY/zyxxGR
lvi4vjEoSmzDMux3IxmO7WGAXDpkUHXqWteCMsYQBmWx3Bv+zkzZgLvtIqHI0GGqnGTQf81nMRz4
UYUEjePp4ai6g9pgbr7Q7HA03NuefyT40+yQU+G5HoDLjG/oZ2kmlmb387ja6ag9u4fTXpPBUtoF
4GDZOzu38y14wTiAGwKm/E3PIMjzjPB2g65p49WjHn5e3wstB26jY/cxg6zIChyJnCHxCmCouOyq
kZ2OLX21RWs9Yr4HKpE/pSmNGrK1wgUh3Rxb/ZbIBZCnocxVc7nbtjpqrNyMJnVhSGrT95O8APPK
I5PaKACxWeKlq14Gjf+zrJQzAZHf3HZn1YECNjo/joM9kYY6Zm7d7DOh8XIvDp+Z6mcnWGWUD685
/letrMT2DpRuMbvGx7/7irBAAZwKTL+8iSRiiJ53Di4JoJO4FXxUyMcKDtvl2ly8CCpcYrGy/xjM
GaTgweV0si8nzqUiDTz006sLIBLuXqDBZ+Th98xVOMoUUmrsw0dvlML8cVEgP7qctxtdaWD2q67C
5zfZciIcFzgQ1NrlTH6btF+tM3XHnQjSra3yFEq6klQs4qv/TSApjlAA4rga3ZWHRPEjhyoDqfOa
0vxnKPAb1vv4hu5bY7k4NR8W9BKnCT7oUfjU7aoB2VIx60poEFHR1C74lCGvkYfSaRzgE1A1um92
xJ1C3xwvtBc/pqUPfWAK2OYX3hAwfzRpyYQ/3+bXifFTIwq5mDK+0Xv7JS3L3jR/b6ktbeD7hyCO
fKFWj07IE77awx6td3II7vqx4nU3cMYD9f1wNq265q1DojvTksA+I9Z/7HQWF7oR9I/EOo4w5CUz
VFkkynJu0m/T3G73ID43PiRuTeVGBionVow+xXK+Cn6W7Ll8P6jw4F7IqXvYSmy3aeaNYNUdyOci
sZV43Qp04BgK1idMASan3cih1enkGJJnHUkh82NbtQoAw8OW2EsAz6IAS9tzVGQbkUcDzY9L1//n
AhswRJYK8+UyRNBsUJG8E9CM2BogcP62XSNVZCHeY3zrEI15y0EOOILaVanRgiBN2WdzsvWw5V6C
0i5Ng19rD6TonLW03mPmasTYEj1ELYcMtTdnIqzF6fqQWxRiJps7WGLri20bwCLRfB9BjZOShnpJ
PcT0igRMfYgKD8FSAY73Y07JqflmARBuwbNTeiqSxBySMlshP2aNQ1Zmo8GaFuw6ohAN1rh1hewT
x6z0nzf+uzSmxZ4GSnuH3kZmQJZZ4nhWBsnR5RjEWS1DEr6barAV18sKDAJgIDisQkNdZ3YVH1Rz
1aiMnza750SjJksvUhh+vYQj88sXctN00ysCvdPij8qOrnDRhJSyrrT7KGrqDsgYBV+Y7kkmcPWP
2FFweV+Ruz7fdhfkF1q8zx+zy8L4G8zHmItCxPauk/RRUG1rqFs4zQbb7NaAhgS/G0Xj34HSW9qV
9BoHYxg2t0ISTDcBOavH96JD6AFiJYeTK2FwJv2g0fT8vzpTvdd4+2vHFdWlJa7WWOPCn0W+Fz9i
+HNH5vGR7sdSeu4lIie2jRqkgRuJWTh2TvFRL7BY5JmF5KsA858z2Tt/i238PA+qKcDLIgTR/s/M
sHvSX8NVm1Ts0+SryI3sHqS7mmHOTSZrWj9RO6rJj+YGKuzKFKdmVkb+j7IrJG4IgOd/JcMzFODn
yjcRYMHr0mk7L6EfuKnK+MDt/6o9GbNHjvlREO7FiTDu3wi6VUf4BtXaQ/nwU/MWAarYZEPhakI5
M4Vp16lKxoF7zOe1OTAdHeEjXY5bivsaoxu5kcnnHvuUL5BTSKWpMKv1lIufRHNctNDom1SRPGNi
QCl7eQDQp0wuDg1WoglWzXtoMmDxvBjCEYamGFmLXrtM4TXwLXKOv+QYry+tHTsWDyfgvuEejxo+
XeZ5lraiWc/NCiTV1aRYfuS2EnLV+KuTP7uYuUMmtLtiz0lhs2NlRrD1tK/MU+gflrysmTLThf9B
rlM00j43zMzkh4yHs+CLqOiIAZYrfDi6QQf/aINV8oeKw0hjl4FokMdXR5gyrFCz9CHBM3kbSm3b
EyO9E0fRYVZerFo4gzYDGwF60I3S/iF+EDZ4Lm9NDPTs4WhRRw3LsDPNBGBCbKQ3F06s5Hw//gLu
Y/2cNM+4Pl2shjsgpcfwKuPbKnoFu7VIrlBUDJhcy0PzhncR85ejjGRwwShdnQ6FP8dmXpNtVKtF
Wsc90MFS2imSfI40iI6h7jyFUsuE4YXj+l7l4IVcXkIYq7JLASKlvvhHzZbJbuPlv0vN4XEpXC+k
2C13iiZsBHCPJtnqotpm41cxqXenBYx7b+hk2jH6s0pkYAimStQABiaxyx7+QgGKIQAra4dlzakR
n2PSgNCLq8yPrUgnAf2DbfyhjjXID2a+D9mMyAJL8SgTi+77Dj6JKTr8hSUeW0SzfgJDNt9URQ8T
DHyDt69wGLxpnTFaMq9H3vnSh1tf2OvFLc7knu+nUgDpjA2uztLJiUw4ceUiGzYrQ/0XHQ8w0T3p
xpHBOrRL+3r1OUajPc6ylqMxgru5uIveu13Vc7HpEb9UOgLNWD7hBx/acgEAj0MKTEGiGfF56NBX
u7VFBSoOaZglAr4XdaDcHJCu722bUtu8tehPh90b456szkI5bJ4PH85rGljBsHcV/lgGxrf3jVNc
khZyM47VJpueHiAnaVfoYdQItNWqCTrQvesbeSpfjigtAOpvb5ALbhYUe9OsmTUoXSUF32zUMZbF
vu4picRym4VglBvHLIH2GkzYhuBP2QJZDr4nb8kZg5gSrxzcMZC00328E7YB2By6geA8RG/W3YmS
72r04MtvvCm7FgY46RrgOPUEZDXnbU5AvoM2wsUC6RnIJTFrHkUMeg1gbDdrrkB+xda5bklClamT
CGNV3X7O1lV9FtKavp5n66ms5P00q1qHedxPiTLjimgUskp3GPZ/HgpOvUJfx4HCQ0x3Ht0mXNry
AXLfZVHZlAnZ+v2SdG11MVjPHEloOpUOOXMVCovh7PPujZ4vLiemw9XTvUgv1qcGiVNFYLRpvvS2
q/gVrFk8VXClUcANFEG0Gh4GhkK532HmxOuRLGOJYSe5LDDaC/mPcoHIMWRfLCcBKnAzhZe+n1u5
gbvgbvqdJPbYGcVp8c6KnWYzAsjZrWUd2kautFUasu37P1IlOm6ruNSpbcoQ1V6TBDdb7dujT3f4
o5401KSpff69Qm830LRSFWRCVKZg4JeKr01d7LNtLeXasHedxco7aFq9oH3hv/dVAnbm7uCAOyew
7DQpyg/pAtGcin9RFxUx9XbB6Pu8y/6GyRjO5WfQjNW4yd3Zu4Ea2MzuDKZFNWb6kWfl7Mu10von
LMdvWpqI+g/IO9AIyv1KkS5CX1QuPJHjfQZFx03RSPjpvhStn3ocG8ZO8uyGfMCmTSWOW0p/NLR5
hwp/wNmtYSQG1y2BQvlAqj7JcRJ9sxGSuqNpy5AE3oW8HbszqXSXhbgX6wXvp5oXqx1l2GI9l8jh
Gzt0YDBOONAcsY9xKZ8gkiW0Cd1SweZVNEICwZgf00PZ7LX95vYS5DX2XXGj6xqhrKF+9KyaOd0b
A7eNw+OD3nX4gz40GmLpmYa0eGN5RmiQCPg5VobOFHMnWMb6DRuEX/5ZQ5OhRzevRt7xPmCSOECY
srPHBAEhUztTp3ooOP1tqkQt9AfP6tqqDI9a02vfsfSSPy+Xvy28FItWwHiaAEv3KBBNd4e5/5Ph
Ufgn7Hs90LjsvKoSoULU+a8bS9miYGo9jrxHsKSfZZ9zG/FutEHM3fbaPedKB7641jFKMhsuoOlN
4Cf4k2oP1U3UeKz6lwEbdX3ZWLWKLzSeFRrdOCohKcsLMNvFEfm9Z6/aFKGEpteV6qk0M/TxL+mj
LsZsDvNzR+/lEZTYgY6+MpaH6I7LfWSL3LjC4UczqZq6wkDP4br1e72I7nyrDqjmuFgEgZi28GCN
Y9v48k5oOfMK6TZfwBMh/TDkbcHKYEHLDzztg//hVhnTyyPYPBw2kUo7PBOQE9fUYrT1OiMzS9i/
tqP1tWNAbMoGSfcWI8jeOW1g4Qz4TXUk0Phrmp1KDS0HPML6CcjFs34MFrP9+7XpHz5AZdVDaK1q
R2u24qw49Vh0b6QBI/zhz9HzJh0pJ8JlhWzRl2Bh8puLBrcAWvwQL7q9EfW6ji8Pt48URM7tCS2C
Ux0Lj1Z+Ss1rAoZiteAK2UI129XzUTjhVlNuilHZpPyHDrlVzafpme3XI9fGdBL2EQimN3Ojo2io
ghlmZlJDkE3wEibj0AUkByMbz75NWOYwTSAzUVOCJHecDVEbLoTclA3dpsqL0uF9M6hwCJm1GekD
etuvEnzrXPmJfAfMvQT1TZTo8N7M3HjFBkDl4gcRRuTwrzu4sXCt1Zz1SlvRI6ZJrmG5qTg7fopn
BGkPCY+I5s4pWUAzy8fZegMH/ZwHBwrCEfX1u1rSo7nDjrw1cpTGJ/4UDRKZW2oxi5YaXFyl4/Os
msNpRjGICOz8AeZKNYhikfGtPTz9WqSLYyGuoUIz/WfVHP4CI9EkNiKswrujz6D6hhgdWuTFC1Is
mNVAdQBYsHa66EKq7VCy8oN8yM6daQQzSrNDcm6yQYunxatrZ9Td4aXBbYNWxo1k8fGvYsZ1Dy/R
0jpjy8kmcZY9rE5RxgUNrS7a8s/EZXUP82wm7w2YNA91eqQ0xgTYJRtT3+sdB2lQAA2VoKllqLtk
SsL+nvHZXlmVuL4TzmyBOdec531ME0B9DBz7e61OTy60mBqRWEnQ+J2tHFlZiDFzpcyDLerYsTJf
F7PrVNwVNjH82+iJXlv/weyrTgUETTVO747mS9ClK49QDf4bhuLBoEetFCcBzzyC3RJcBnOscb7l
3qE2mUFpcsiupB67bIsPSW4p+A0k8rT9e2dQL90Pcdt7BED+C0zCuDfc6RuORSpqEHRJrubSy1Yq
oFe7YT1dTMLoXnOy1V1tEC+Zzy6b165ayq4ww2UnMT4smi3aC7mIys+RShQv2lZVVzkXNNmDbgO2
4+RK6Yt196RPl1o0ehG+c/qjpMeNiYJkscXo6YkfxPVHTIonV3rKt99KxM8GcEteJaBuW+65Y8qP
sZ0YJelXq3Rtbbv0QL0ryYAUKKiGuuL8NGHAj1Iy1cTl6rq6lDa3N7UwUBFab/WUfNoJPRMEfBJR
wytgQhabxHhaUcYPcMeFtBgwigb8ukFVidAwpi0Or7GcNGVQmDMn2kEhcsucLO1lI+9DY5qPF7Xj
ucpqpDWHkTQ+XSs4yiKz4Gc+5tog20EtE+OecHftlym2zhUsOoICXtMxaj5WbJl6W/KaV9vLNb12
tkTsgftV2hNIjxv7sld2lxt23eCuH9UMcfiUEDoNN7b+GB5tI/boyl1sVftiJ9cbcCy9fMIfaIBG
M2zBaVF1NhtgUALB+xYjbZ7rOFoVDxq/XY0bVkLYkvSGQU1Z5XzCQKjlokxHmL6n2EAd6SgK4PE5
mxbeCaxniYLX8w3PArwT3AfQnscY3Cn1kcHP/65yLZUfnoOHJv2kVTGGZ864n2/jcGODCCkYpkAC
OQ9SujdZpasurwY5w7lNCmzz3R47gtnuFpe8CLRsfrXJOnUGg6ecmuMf1eRFHYlqmY1ndf77KqEY
Z5ppwUFHzTV2iZHSUuhiBt1suPvIrOGKdakE/XREwnhV+y0zHCX6uebwEZcSiUvhB1hawzRGJ5iV
EtLDS+SqoaVcGpOqcIN+J+9JsGxfP9OTbCf4ovjMIrAa9WamE4hmkyeRiLR05TCXu5+vqYDr1O6t
oBPxidRRqjWNq5PQA6tPS2/upDoEdOeBkkdKphYl1hEW5Y+LIrBw59k6B++U0NIhNJ8pWLx5Et4k
zAue76xN61b9CdoS4n/FA8wu3Jx+W35yO11ZuNOS8OLslRfU6NGvSEKDihQEz9q8W9/+RDVIjz5y
svjU90s+gw3k1WTAm8AGQGYBTNEODuzJSZQBMK+kRZcLiGlEFUlqmDmDcgUqoiTl1DD90HaBq0cx
OuvIyVZiaOx4Tmua63BmboIbMfWLYwv5PDvvlH6FXv4Ia5FlBCs2XKngid+mqaOqKNUZaX/58pf0
jijuw8qjIdt47041lXHO773KXs/i+iKzzB7Mlaw0fRpbcVHXc43jn6/S0yq3PTGzUv/DCZH2pkWp
qQyqN9DSUlq+Yy9W4bTo7+RX11jEzCv76ob7pntWo5Q3FO+BciX5JsjCmJqydJbvyrDQ0TNzwi/t
ywIIDcFh/1DnVarE1PDPIjAcJkM98YHhYmfoHgp/svKWvJOBDIb4GlI7T17b1iqFzfNxCQwsaBU9
lv0ejHWI/renyoC/s7TphzZVjvqL5OF/twgdtI5G6wHz1eAvJQUB+cetvaMavPZhI7GEUyhgaSdy
ZRuQui2TGZYuDIu5n2kH58c0XQ1zTNEqgablvSvB31gvXx7JcFmt/ok0r0OGbrn+zwzkL4PeMqtc
HBsvyM4X2MPy2Xuzgm/MUoYA+VW9bEdonWFdul759Uj9zNRgCrqKcJnFHsXUjQkesxfvHR2a8VWH
zfNRlWdcI5nevqsjFQE8CkWB2oszVSb+5t8cq1SxCSPUxmXdnibK8zCyXs48eCg9LC3x01iXObRv
7lSuaFgva21gDs6JKNWU6nr4P6OwdBwwfbRoK6c9KtvUjKDnWu2I/IRFiECMuAM2b4cNK/E1eh1l
W/ydzwOD2OQ55q+T7vnyZTDwjIMWPnLgsQytpO7AmKlAPhFT2mY72FQ9HtG67ZhGROlknWSIHcy5
eHPXZsomxqj+iIkuyNZlpG8NvQroOi+s4tkqZCQnviAQIfUW4RF1cTnzNYdOX5t84b9mGUGcQE4K
OPSGqtNHk1dEXZsCvNXJnsXekUvY2Bdcj4Um6sO4cWQFyvkxFZNGIO+m+mAJpbJZzV5FxR3wpH8x
O8/oKErvfLdurPV/Q5ZrZyCktTc8gy+9IdB3kq3CmedykYUbU3ExxXKsVzVWVdiLGd0QL94rKwJX
oP81Tt21fuMNXAcJslYUoyoRb/ExiEbcNAPzUKL9oIYScu81/8UZX0fgUP+m5omVPJ//wN80wNhQ
A2nY4LNew7yM9lk/b1q2As5JPtO754YWg5vsftkITmKqTf61AkwMscrvDeGoHFODKJlXYJqRMTV+
0mf34tKU43+QGcNKhMwIQqBsblK6wYOA7mZefK0KxcOeuDuOZvtdyN+u9Lac0ebmlx8TrLjPlS/6
yPJ9As8SvFGukocBlLBB9Gmgr4/D7UOuuPJXo7T/cVnn4k4nzQLAxnlk8BagihWJBPkMVUBfJWnz
u0TFn4hHSBZ6k+qrWu5JoD/+HNlu5ryxDXH+W8tG3A4uuME/DOf5GzSwkXKvSlsoVXo0k+3jKlHl
dW8gGJvKgJ/CvUhssyI8rUyJQhA/J0RgwueowdN9M/smlBIV/wUB/LODU70aIgJSEfw86E3HFEtL
QZhwDwDRRBDLchR8fWt9EGsg/3hgc+cxe+BYpB4iETt9sdcjva37bKpfNfrsv/0dAv0BaA7tNj9X
ULrFLtq9c/W8sngKF1F9/nj2LNRSajhN0ZAxc/3qXD4AVUWhHn3bW577PWcnqBwy8RGrcHVATNdp
bAoCXX8qKbRJaxYk0pqQWELcpfmu6ml1urr8ad7qtRZWp5sOQgbZrQ4XUJeUuQlH9siUVtTguAsG
pxvJxntojtXresqKbM5p51JQMGm9KbxUzzrVSGXGjSnA75EEyyvgASULOPu+BdP/RAYmKsvhXlUX
79xTlTeayfZqBk0ptebUfhWSc1Q+VVdu+PIo7PD+unloeSbHuiupbC7RboEqFvY3+vXORQn1ZGCM
gUFDGNIpvwYBApjbSbtUSVMOdkYqyYuxZEekjG9r2a1O3IdL808QoocHha3M4EuEIkGrAMIFmEsF
3ajTE7JJY2fF+YYI11EI0RJPAJv6YoMvRi6AvzONU/VbLgEQk0tIZx2NTDy+B4y8Nb0UKscHY9Ok
QrzjCnRS1KH+3VEz1IzaRRbJJ6+i1xQjHXe0uxk4Sm+KWC4n4yrkZQ8Lc0BVZ4by36gVudRBsvU6
AeracYFQPKEy4Lt4lpd/cHAiUkcYjOMdQ/XXkzHAjadyRgHDWd/FIOd9iYPS0lyshJT1sBVcfnJi
YM8LKN/4WvMiFkA+nHTa5ePYltxgvKeoek6JuPwDc+KwZxhFq60aLNfUP/79VFW4QUlq6gsz1bkZ
ViwGu4R9xdxKrkH9HzN97LFE6rvgbPlpnd+18YMwEeNtIJHIExDc+oq1d2F3fzaD81qlWmTG/Oqn
fGkiMu7ju2eET0xhs/uPzwJML17p4SbPEGklACCQcaMskgyvDoJUhNtplCUWvuhtnE2b/ihdSXeO
i78bReGqauUfZBYpM0GTDfA2NE9Dd45Q6PEbE5iFbgPQW3VsVYVsYGPyoMtpVtmqt/jWUiNXtjpk
hnu4cll3PM8ijQUIosAJYg06eLJ6zKMT25cl2dFiLnGd/9f/HzFRlWxV6xmnbgKzsQ8maL2ODZZP
oeSdzCnlW9BeNkE2rj9EtB8bBXBLRyxTp4YYad3M5kA2O/kAlnP+LM1jvvflcGfFhkuTHuaamk+K
JPyK0jn6ZJhbbnu0FQ4bUFhcM3jAXXDoh3hEMhg34ig2r9sxIrYek6tUGT3s+/W90wSqjWVtqJNK
QjKdRU1QdLB38UkLcg9kWKkQ5kGFlXvfIkveXQ4CbDDI5yvWq3yqn6bXvUea3YMJLvBTcEfqvhhy
Q9GrSLc2IFGICr4yqYwrAgdAFdjdXxuFmYQXuCTLqIPpgjqnMv6S5WC+eKeKz94C/tuiaAJdzl0y
X9v4SY50L8cMLBQMHgr71SWTB85xySxo5ltIUv5VQOK9GChmPhmZ7Gc09gYKIcEwjEd7NgrQ7r0r
W2CR5uZ0HClFPwA+6+c/+L6/OqGj1CXyvrZAttYN8D62JoZ80jS3P+HlcL09/h7bDvW6B+fkbdMY
ew6xjFO3QiBp4u8L7FL2LkXmObDr7OO/YFZrJ+BUlayWtp+eM3Mr3/TiUFSkXq5xKQrG5qfvl35u
a5xJnUbDXc+xgA133aFAbAuGMsTVpee8UWcWS58rPFU1DVnluIZuyo8JbfwcwBNgLieGQBqeZVnd
wcWzH7Ya83aQ+H7yxRjFk11giNSrpCgtZPVl8NNTY0VvHBrqNMPNVYnV9MEiU8jg3N7JJ9nJIuo/
6RedCS6HPuLTiwqWzy29+O0TD7PPexmrqC2vADvPl9bmZCWiMIpsleSY5tc+od4JhU74qj+oUs61
6ulSWCiHuvwgpW2XSmEoAosjeGR1+1/whe6u3LGk8PP7LWSBxUWJoIol/oMpFv0zG24sOxrPdPc4
szwzyGF5yItXtC2ApdIwipsddeFbCf638sZIWogHX1kuVAig2SKA0ZaCiFnj6CCPKiv44uCUzZux
QG0tISjp0Uf2qyEN3yWRqcQcajJN7Xk5f5JVcKzG1LdezmRRfGeoqbM/MlJT+credkV1QD6BzhKC
FzwvL7huKQJ0DcnuLtnRJWg+E8afn3PqO0QkKnmkhhvH90dckk++DwJ8/SdtSmQ40Tk601SkimhF
hgAvkKbNWqt6wmFGwU1TXA/VChfx5qZfz0tqMmgwjWSgNTZ4x538keu/79acjfLOr2kH5JlmGU+M
/6ZWrSuNwBnbfGlYsL3aKxaB/6TeWPuxmz+WfkdNcl+gVbLsJ6VnkzeGul1VG3KzOq2mkHCy557O
j9btUudt4V+UzkLo5R4lnJRSM3CsEFWZcGQTKOiOU85ojmiKDOIKN59T6EdkMHA56pzfgNw7uAmG
UHccgf65p4+WbgIhGz0W/IMKDUGsGdEnkr2HmGRMkFQlnpy2ucyFRy/wv8ZQVSuK5rMw/ZZ/1gtb
un2JDSfuYySqMSlJMOdrBET+xuUdjg5NI4cdLcbAX3Q5IZqUcIrgC40OPA5OsXnYw6lN4rj6jjUx
bPD8LhQBxJmCbwR310JgmFSNeSxkP/l8ImkgcUNEtdnLWij046pKXX9X3UmTWMLt27M7k1a+SfBf
e90tz23uNo8mZU30iTvb/NYTlUHjP6FlEirsVPIutmqBkrt7n4XWhZ48yRRKxxohoXY2vvoezJCP
wJ36Kdvf6xwunEFvtkf6+scWXGSEiLX0lKl4/vjrmAXEaZVJ1Bp29D/6Codcq9Sn0oMX2aEv2Z19
89u7jL3pb0sQIjPSQ9IoDFyVUzRMXpk5CzSELnYyYdkfGKoyJDARLW9gZ6D/cyYjTSgOplG+nCU8
0olIrQXnw8Hr3JaMVjW1n7woNbYAjLYasrwJ6VmEbstfiWvTZV6GWDyNTOjVfLsUc14IcORdLZOY
vQqqqrgy+dQpoR5ba0oXk9F01vnZ7TUtA0+DyKLpfRg/6CwV+Qmxv3ilm5wQ84/25dB5iUIcm4Hi
F1S+qbntEFwlIccHgTDkQvnIBi+9mwCEu0UArGynB0CBR6w65mA3YWnuTbPCHNcBtV9IxpW6jnWV
XDV/6yIqTSsoPBOIyFPcq1MBK8hK8EsrL0F8EGIZRpYD7jcnqvnKJXquPibHB5BvKgcAnxBjNVqv
iLL8qGoGmkOweFt+La2abn2EA8vInxXzO0j06V1hCb6zEqpAjPkN+nJEn8kUvD6Btts8Wlfk6mll
yF7OqOTHUCFO6Spuqf1NNXVJJeJEe+YgmN3/Ymnh1MFvG8ZX6/weop+WWpNejhZrtalOtj2KR4Fp
4MMOl+bPjEWWpOnUJuZtsqDqeoZz8Qh6qOekBqq1aX/2fpGruPKtu+qm4MRgMRj1zeOR0K8KRtjj
zoptI1blnNgRM9g9LnaJUu20L4X67hqp3E4gOwjR1J3VijjIt49MoqgA+C6Q5VV8zw9svoeIrc70
dNqAotuXsRwoSsB/QoSZfXlCTuNEm6huDP2s2DoHUS2EV7dhg2VN0vSTzsS+VvKTm1b0QK+kFej3
HALd6a/wiX+XpVFwM/RK5vuL8bbbvwFT29GzL3+C9PM7mA6pls60a1SvlpfbZKCUQrua2HR8SaFs
k37x1qqS8F2BEgqX3tHoW6Efg/5tPDh+oCGL4Ac0RTlkhMcR1QhZHYphmuRREfBqMHmFvoYiDhCP
DW24wK+AKbCkxv+u+g3QoOi460D1sLqUfARakYPEoIEbuObR+10kgtCIuJuWHm5yjMT5IyYJUZX5
tglhzibdRFai9oyCcUYO/yGyOdCLZHrtr0lKTfg0VwZBJ+voDMNevnCAa/0iRVe/O6dxeqE+mqqf
5cqC3ydBKHSHWxiZbELCu+Yw0NGwXmrbvqfnBOWu1IfiSsBtKJf0jwKfp7gfoUXnkLITpvGniEhb
LwmUli9JxRN3ajy2aID3LtG2Y0gWF8IN8lTXTh20yEK15xOYMXLSK29HOW6+D5d5xD4jOLPb7dj/
3GulQHBSqa2DotyRy/jH5yIvg+nfli4/ksy+3nXW8wNkB2cL2WsMgfFXtcJJlHvHaXuSko9RXB+u
36r2lN7NsRnw9Tr9XLuOxykcjeSASWM5lPqCyp0lWfDjlFlJq7hEU4zq9Vu70AnG6sSEuALOOpem
3zkwoq9VXVNDBhs1nh+HLY1xWhOxO4Crf9M9thGbWxeKh1/G6yet4fOVTC75nWdNpsfxXU+me3DP
ZVAQd3Mb/AssqfHzZk38HQBevJ6csJOGv+/zSPDQUjZ/BUZKl4K1zlHMtoK9Q2NiROo7Iw3sjjRq
w7W8Qyq2ZG7XQfAwFVEQZClNPM30AcqHr4b/dBXWPpNLolMQQq2yZWesCMS8mb3PN1ZSk6d8soOf
mFdc6dRtY7LWmQ7ziUmUX6DPykFPkYSYC3n+gZS8GkNNxJ7PyaS2ErONRBoLxBb3Dabbvo/Clsg2
maAIHc8ezIYUuCuZotJZw4LTWu2pY1kAVHqYTdi5ydiKSqgfKUxaQPAxkfpEnHcym+/CrP/1TdPy
9sIt+vb0/RZ1ykfIbxf/wFPQlcAeGbcdknZqMAYCVj2c2UYzpANFncLezWHvQ9XTueOtGeJHyeNG
VWJrZy/jKSDiwutlvscpCARA8Glvwtkm69ozMQVFDkxw675nikIYUY5+nfzIb8sxrPEmdTvOz5/A
pKIWk9MRo3kkR4cF2eH2+wzsLx9Bqggor+QQH18FH4I+2JZH+xsRkA/5PfM/RIdxDDv28ssHY/9D
NmHukE7lyPes5SP93lat6c2GLuslZD+oTpFB7HoMhCrsf1Ob+De0AySJG67X1Q9tFXB20B4sVmIL
u3igjotH+Wzi0Dh0c73D8LFCjVvZ0Y4bEtBtNutGKB9PU+G2QkAUf20QLFcoHAbcZjm3w5O4M1I2
Bt56Us9DIBhW+2aVPdAiZqhGWP4JzzWKV7VeFSwdFIfQ7uipjmRjhI8TE10PdTb8bScYnjOry5+y
1eESozmvOOP9mwtjJ3CgoyAhuf1C44DaZzkZo+NIrUR80GSTh90lvTuqZFbdJO8XkmDg1+JFaf0I
Wa/fRioK9jXTAlGvw5wQUgtqnti0gSu0g5dFshFoBBinLvmYCzpizA4c+UqBHANQq22gm5BdAE4b
V0FdQixP6zw5QywJDh+dbyE39YttUYwxAktyag0HCXQjdU67rxAjlQb0GaIVM62timkjIW+Z/mJT
iOYZ7rU0j62khPvXV/1u/ETKJ4XCuHbCbGOcs8f3NLkiUcF3+otDdFl+8IbOe9/ZY0olEdOigfLW
T7QUWT7tUNgviwTVHtbnkzyXR3XIKomcD/W9dGCY8JhuDPqJp24RmZD0GcKvidiFURV1e23k0sQ3
qA0JDLxyAD0BAwWCxKnCN2+kYkn/AJdTfLHf9wkcs78pCijmPj+BLwm2e47dwETFQAw74nHF1rWK
B50OWPsUbJn6EgxjqsPo/PfjY1lW8Ojn/fUmYn5OpG31S0X78c99SiyVnw5QgEA6NDB9gczgnvLy
U3Z8gy4jE0VZfLEBCN7ufk+E38fHKTwcG/pufZDFZ4/6k+z5c1bFQ0rxImg4pBLe+YWJkMR37IeY
DkvzLpDdU7nNoel9+MapkR8lsxYg1jSufNs3kLPtcwwATggG1BBTYp6PhdAdlX/JFTeig0qGQkp2
PUfAvdT5i4WHFWPvXIVDRN/2OYtJZzj1MA7n283xnjQs8sX+sWZuw4u+o1fWKDCbMsY4KwxSNK7f
S1wGEa0s2T7buk9CU7KC05YvGsoD9kLoFg4W9A/NRB02jdZk52VLJ/ypokxoV89VvWYiZ3so682S
c0wwJjS8n9JbjTxXiTToT4ASlri2alSdSCqoHb7iqj8/QjTys/i143MXVRKfPW4gzxHRvdIyYBiD
7yzt1YcCHLtqNDHij3JuFMD3S8FEFBha0WRocGbAIIXdzudmyqbu26T0k4gJ+p0jQQ4+jz6btoid
l/twKWuV5isissMcbGVwIxDM4RE/jQZOT1oO/YX38tnoNEqJGdPAOFZeV7Hye23SP8F/VeO26Wop
rZazotTVlivDX1VmTi7Gh1DXV48+IonwCzJslgKFcsnSIVMg5J/O4Bf+92Qg8vkayQKGQ2jfCFS7
Lb7Z0B4l9pOJMpKZnen93Gag8jGxHhQ4hbVP18U3TqZti+xkCNK38VB1z1lvNUynWXdv/9O7n6PK
51PP0Bh0VAB76mjSpLjCUuLRAWcS7dyVts+D8rI/Dmn+qHXbH+MMhZNdxUfGeCSiRJSkPt+Vn6Ft
XV9cVcFv7eZGLWfH4dPw9YQDcn8UlzMj9+P8pEBx0GRjfVssEnrbmlvhAnPG9bokKct4DUI/wqw5
jTZ1oG0Yth1VEbzHgSGrW9AY+k1if0vmwQbe0hMCv9U3X9SCrSh+/yhdv5Bvt+S7IwwJ3dC4RdHu
k6xMaha+y9UGiJ/exjKv3pB+pQXea93FhOIK5318Wd+enHK43IQqn8UpX4YH+Nsmp2Jfmm+i+y+0
JnpVgLjWvFq5qHAugCtc7xDWwz4U2Duxrom2YpMOGFwZWaCn0zDo2KTKxe6/l/pQB9z3rVlaT13G
sTRH8t7gCHkUeYNULK4GFdVPxWU1NroGgB7SYQBYLQHtPu6CLUUsgbVDQffEk9f3kYULGke3llM7
segpM7ITrlXi6bPi0qTiJ+3mPPQEHYgQUvdpY11btiP1JHe6tvMGhbOdroJErIU7q7ctQ3+NX2LE
kirQj1VRFFViuINe6+2+Z2xfTwd4sVXCPZDxR9hPVeadzBShWMKCiAhN+Fg1iPUS+KkrOIprBWSU
hIuWvkop4p8gmVfiosH9gC776piaEfAlOYvOSjW6dmUO7YtmH4tFKC7iqK1tH5eduCQEWSzgN2/b
KNea4i1T3w2NYFyhNsqVHB3dPaYS4N97ir7lW7BCwiZYaZN/xolWLOPJesPhwr9hFyIeHiNhLyvm
Rn4lfLQAeUZx0H2iVYsnLl0zkH8xr/6cg7wxC62hyLl1CXB4UwVEL8Wxhj3OPDz4nAriutrm9lZ+
T56mgYMXEXnH5lVJGe8rj7Fs39omHcPXvh0/1ujJtUqIyc3T5p6SNB43TuSiZk40GULZSbpA+wux
+8qiwpMddsyQaTAWLSvgYmSMQi58BhVnqnpeEvx004DYVgB5+mI0xRP8sREOzUoC8eefApyLNU4K
JyJG//uct4nUlTDWekFyoMaZtgeuOZL4HzDSciBYT40V5rhV75ZJooQ6INFqEJaEO3wcP9eKAMsf
7l9O80LsXirtRr7GxuZpJZMbvTvtZwZbvUbyTTToUIiPgp82MSREYvAHEiAadDrSlt9ed/UsjtaU
jZHQ4X4bSIVbSsNr2sFpf5kuY1Jp5VGL+pCZ3zoIhuLw8k5j2dvHffulgrodYroQp/AkDBTjZJDA
8kVt97Hi9H3JP7BJNVNE+3uv+4ai7LxJE1LZk80Rex1t07pVVJn2HS60vClL20cjuKEmdbfzWWhC
LYYJTWyIX66gaJSHUdCUVjVEnkrxE3MnCVDr04+T6DbFFfKbQ5Lji4GP050NtvvnmbYBMIcyf0pu
1PkTC/kxCpDEgGY/uNuU9S9gCuaGZNfiQLHHxg4q5cxA6NWnJHkCbc1MQ8PHBWYsL2xAOQ7raYew
VpVGVSVu8TmgAxdnGINgRdE6da/BHYr5goeTZ9a0owpzdpjU0ZjjUtWlV/sVmeHRqEFSJ9yREKkJ
SnevbEF+1wyb2xuXcTBHxsDUTvnaGA1GWM59mxG+loSnBdt5/GoI2C5w2wvWz+H9y5OgBFg6CMpL
WC1x7vE9LrolZPtsxM/dBMt3y42TThPdW0ZlesIsMkDrxnjrkmW1PmsrGI0JOCOQ3AiN8ED9snSV
NsKxQyQRwQr7cJ6pFRQ0f7QanMVo5h3oKex1wAkiEADYCTPal04susqUpHKpsC74FkvcInY/MdZq
jSTZcbUo0AilA3S5kHNilSumsEij48Nsts/XFcnHhlEPnla1km8NPentS0uvPfiMIGJYb5FLSs+d
FKrMUga7g765RLOQJwp7wYHA5d26kuBrb9xeJwPCAnlKOggZTyJjPdxOd+6NFGkERc6xz3hjKUWB
F3Y/FkgXEAGmwvtO2+cNO/UDtmmFX8gWMdE4T6faxs2vNxOm9pbE4Ndj+PXAxEwQ/4euEE698Fwr
0K3EUPrkeee0ZMGw1qnuSCCT4BqtcfJ51IsFdx/yO7OLZxGps901KmOkbk6rNccOabtKdnvJ+ERN
hAfRqbsXa9coL7BtHOZhMmOiYRx3wd3I50zmKIKUDmDA1e19eSFmaL9yn+6LgY7WA+fV/MseS6P8
yD67ugz2JtoYJxophCsMaZKKscNVxrh/7apWQcpfqXNu4fhek83uWSj0v6iLamA+81qs9ORXwWl6
PnnlwyrEjIW40rEVBjlLdYT4mpHFuXGD747HM7kkw7/iBd7BMx9fr66PLXtGwutyB4VKF8F+1X6T
V+E6QaCwEb++Dq54UiKv19AGx9LjsV0JRy42+2etfSEmmkLR3F96rxz8J8ArN5X+9gM49/qlaQlG
f6I63g8eXqQQlVmBhx4GOkRo/5mn4nYbSNOPjpiKBedZxJ7BOI/FQX77Bnd+nbCdOpXDegJa25i/
ludWzN10+2QP5yrZ70lm4TVJkMrqOg5c10P83pn3fJJmIqtdxDtkQJ1x8FcyxuSChNPnvOCBtxat
Whlc1G/Kkb1KEzYZ1orHsdmNETIy6oek1NabSY1xJr5m1hyf0YTJNHcUPp1g1oCx9BH5z9huDrLv
L03uu2L6J9a7uNythazbvq/4NEoMlZ+J5W7pKxCqzKsRkCGiHY3P5pW8yGv8paJTg9/47buU0Iyo
THM/8Tm4ubQcQjws3R5ap9ZoGN47Henx1gq4Ojy5ZPmRBLwY7rTG+bgCp72+m9REpVcFF6cItzd+
HAHyfBv9tADNxbR1cBIa3B5FpQACXdDmO7jTchd6a0dlQJ/1byIHCztLytOvGeS1M/vKvbuole9G
UgpRhiTWbr/vO1lPac3lzxemU/XTVHAFR6kIL4OAM/gOZQ2y6Miuac8eIynQqGO+rs9NL63X5WgC
VaUslbyYQaU1DVbSzPJAFKLP/ayVcTbpdtpaSW1tkVZrICfUeSvrmwEZQXSh7fCAjvdkzSjmBXwe
HGfjmMJTk0bfFzqGuOYnmp9rwglEO8+F8AMJC86T5Z631vkaTaybwXFEVVWwqeFpe6fKllUfWnDu
1M8gcgat408f03AWl2nIQ13x3HfE1XIFsBgt9aQcYvUn8/kpSDaHNMGv06n6l5YeU5kvnLvwgyRO
hYGfJlZaf5Rq1U1VEFRAHjimYyJblNGm4paMEvcNSmYiLl65t9PQ8QQZFtw7H81bAaFLrqvN6xSt
8ie2WHO7FdoJgS1aXmXqgCWc5WrNEj66RitcoLRGy7++n7dFJPUVvlLt9Hm0v1kbR5s9npEr+8k/
qKswBpCFsDvIkkiVN/ryqjUvqElbeOrtQK9Xn7vwONdhn1tkdMnoJWYMJaXqo80udzgT3LnKrcXQ
ytKdawJTVQtaVQC2CDn/2gbYqnXYQDKK6ykWXlnEYXS5JFZ+xLPQKTs82GgCFLGbGoSN/tjbD+FR
vwXaCzp3BQM4109+mDy6y/6rTWBr+DecAzpsrMBxvrYhUVn2LG5ku00xmmzMp+8Ayt251qOU70M5
k7R+TXwX+tACiJ7bMx+tvuXTMgIUxLsEDhvx0ae7bLRUpvBfbdYzWg5q8Ih7y/pobIWnFc4f0AY3
gWFdShtG9Ncvo5XacjyLw3mkiofjjjwd2FMqdkJNV8xLpMgyrXIKukaBD50EY+oDacD4YrJUlNXS
+dCPcW2j6qEileERDlXaho26fBhoBEba7zx0ZshME4ZAEy4PuXxvity9+g9Owq+1q2+e6dKz+Hl/
7J0ObueWfAxDZ/YL8LCOtPdFd101+nFofIRQbzfxTzBV7Syl4lQWxlWiL6xCFOHCG0UzG+4Mc9bV
wIbEq+oh4/tbgBjCG6lN2rXeD7ZfgGOx7C+0BjWTKmoUn4oHtXEVVdZinX9XKkrM3ka+TW35agCw
4X3xgs6CJdldM4c52nVGdqerf9IutdO66PTGzdSLeT6KmqCs4/CU5g7tsI9bF/beAQgy9I9Mg5fw
ZJC469/Fev2zMCBdyDS4S2GQIEyynXJ+grnt67W71kzVAy/5imZFVYQoY5b27vz5yS47wMMsSY7g
VWDpQl48cdbASwBWPtEd2GCAc/YQDMTRUvZfEEHVU9bNg5BC/9Ju3Ob/Ig6siMoR166+iQuetrH0
GgGVCsVoOWGiL82HX4iIytLsTYzDqv5UHJUfxpuepImuQ78x4Posr2Gow67M8XHF7uTGidSNPUwj
YUZnMSqzuwYHXLEotXxz0BkcMh+m2EZsCtGaReQA9yFUNQnP+ODmUnxlYCkSHMBYJIUG1W9D6Ug0
tqceVP+w0iNfHCvxlKZT4Ma194F+FQEhq/lImbMlyoNiAbfuBQeFy3ynCkVnK9NTv1rHwkDIlbLn
a2uzKKsnSVIgs0EGBdY7NC8z/qZfjVgXIQcSLedZbyExG/+bbAxNiJ44+zxoCAf3NDzK6quAZMwW
gMRo8K0zsvVPU5HWRPoP57nF8olRGVD2JACUo2pCIC7t/JEMCce46D/rUuIq/1sgDTGTsAwWNKD9
UPh6yXKmdmOO6Dtw3vhBIWsi3eZnWEVpmlJCWymSHMZ68EXcKBxo/V8AfrGQPyPXm76nCMc1L2Rs
USvtUw0YMV+N949h8lhf7apmrOm5iLV0R0B6S5rkiwzJot322uVAs5ia4o2wQmBYSKdSEGjYKR1w
/h+ijsuexaIJO7eKmoK+vNlTLpeN7DkuScnAz1doKp8LsWoWr5fQelwxWXu1J4KiVX99NOeu57h3
HxiEpGn1H0EtUpq7yK0PDsTSwKadLZcbCZfjPgwDM68nZ2rRKO7olZLRqUuCoe92Z8EnBvb4QonJ
0ErTRWStvujYetlWgO8SJGuY7Oa/WnjrDDVhaR+WBbGAGRvBimVgy7GGnMH04B2UpjNX1G4NUhe3
VeljKDIIVLVl6LO32DgR7wS8HMJ16T6KQYkS9WZR6YL9HFAl7+p+tsjZM5MbHqQtWQA321LUBBMg
o6PPPRR8Xsu2mkWsH7Gt8pWnAL4HH51sx/JUtGcvs0H4LdOE/LewyK9TGeDw4y2ahn54hIKdp7V7
86gxNMtL9MUc0cCk6ktNLg+l76ex9HUXJv3THs7Qd6XUXZHnYUI55lb83m+ucqJAX+ubqwMsMsq2
8bcA1vOMuzyehqTKROz9/Pe+qdjqhb/E3C8PmKH+Bd8gP3/wmRWh7beQ4f0rxkuJ0jfBJ4Z0iUsV
NIKRPw+7krC3Mnt0JVGpOG698f2frrpP1YfiMHoGlzelmJbCOHOGaeFl4Ly5dUMA6rlhXLj/hSSn
X32ZkjEnB9WY6JRyv6c7kYBlXagV9qYwwFWs44LfwqfRchEYtg4an3jBvtRQnICp8kF+xkK3FepL
sWEN/jVs+FeB6kDIhReXFymYBIn1qMG0f+ACjLoWioLqFx3LHKaGAuK4hiQMLqAX5XjvcjqnWrvJ
uXA+vMeONPDSd2cDvY0Ju2YCV+mcgTs+bhtjveE2oE09gv3bDkcOWdc+c740BMoiSovmbUHQd1tK
zS7j+CBxucKZ+WS8SVPNIkl+fyB9Kb47/zt7o58VRwqN37ry0mbFYGARFmXHec9cBktfScS1L8AO
MoGpm3pKUEkP7hJf1quzNJSY5hO8w2yla0Tzd4bAPrF6eRqVc+E3UbTayBamNU2EGcGf/ofJVDq3
u5ZT9M6ywDi+DXs1YeFML0Zs6aBQwWvJLJ1E/oj0iXQNrBnZuW4eHZDHQeikMxztfXkRTrEHK+PQ
+aBCTAWVPFbF+frsWm+G5knLZqRtdpjML+6Iz1TDHLYp+MuQLawk96xe2inama3QRF27M8+pZf5r
ZeoBe5sJ869KdgC+f2Ye5ZH8hLkslk0cOA+fIexk1KmoJN3BfRNvrF5G6o9vP5yHXNLHTYyALObe
00SC7A5tCljcD5Q2QxQhrxgn1NFWhEUZT0iVkMrW1zf5p+Mi2SkwXUXgnaS34hkrhrLHPzVAmrOp
xtv/JCsSkuOsofKl33iVkb+RjuiBLKMrXC20b5MyVW+9kTCZnUYfqxfOh33m2F/F7U0DXLFm85fv
NlCRLpMRIloV2Is8PoJfSp0B9xyEWKNJw9WIA8dQoL7E0ws2ohB1N4vSUeTT2kB0M+39XNRc4Mh8
Boyo9a772TcQUq+oWRgkh2cV9+C13nqFKZ1McNatPZXO+w5kdiF39e2tKShE/8JbjXWYbjA/GCAQ
zWdX/JE0uy9k+LF9jX+1582kV2zGT+kQ73pFppOSo0JEHzauUfv9X46hbyE7lQ5DvG1Up7NeUw67
9PHx8ecQZRAufpulNZPLit5ZuT6EEizuB16/sTEeMn7RDTT5yb0dpbfbv/6bY58tpHA1hs+LwifQ
9RPi76ek5982Zi5+m0EFIGGYyCMlCCDn0gEZMCvoe7CxU4W94KH5ilOGhY9sWX5c9QEdEvJSpo6+
WU0NqkhfxRkY5tESbkqNoaRHU62PssI2Og4bkFsG54sD05Q3lt2a1h016mLF7/3ZmFehdGzmvWzB
nvoABhWCCEXr1kRtXzeztNxy954K900O7gCMQGtVrgQlPiSm+BeJX8uBKEtVk7SaijGT/k7DWXRq
6UPoOrKQZENb/UFa6EKiLIzUCjbTpJkGao9M2J3sDW5VZHKH4ZMQ4Trh7LBZnRPzDpSaaeNeEKZS
7REBUfUtAdqb78hRaEfrzPHpPapqbhmpjnqF3jKPEAVkM7cDnkIfEQb/bSup64dDMxsDoVONxcyM
SlQvTlKFgj9D/xw4meot6GkFt+STv1ZAMMRrms6hU92vwN6l1q+JZm9p7WQ3bO/OMgvT7a0X0cfL
sH9gJlwtkBwzcpku9YvklXkV3J7K3PntXxpX1UhLsu0KUmMvaREGazese/tKpNP8qjRXsh0EHqPP
LmSSNotfQ312gAmjnqIuiuFJ3dLkxZpx62D6I1X49muduZbDIhSPhDWSJJXqyPdD9jMHlUfkTYB6
gJKhLJYe0tNKPrJcA51M/h8G9QkWfDqob1l+FKx+vAJNBCdNHyjpkPSIjpztHKsyZaqfMEzCpl/B
VvYOVIFY8d4GSFlGEqFkhVBV+fs2VahAyb8tG9npKso1wqcquNge6DjKbqGBKYId4hOKp7oDbx1D
M8lxwWaYrlxe1tFEVsPa8VQeSaYRlatW5/+FZ6wco7DEaWKcU8oF22FbbyAf1/+kuw8DWk7BaLIl
A95sHeU9bmiHvoFvB6owwLYVuNs2XsyoNSbN3VzTtFcIctlVoEGZjhMC+36M+8DPMZJj5BfYUFIj
T9v6lshZaHGWnPRAZrkJpOZKVQK/rbmiZyrLda9mVlBamPQ+SKNkCu4A8ZVnOZo53auyKsJWSUIc
TNUbpMt9rpWt9zPa7KbL1MuY2StG13JTKEd+UhatumTtcq1dac6UfgGVHgZgpAtEyfhQ22sD7vLM
Wz9ZXeHbBHJ+h8ei1vrL0FejmI2p6IEiHzMvu0GUIfSRrQMllHT0lwlSx7JXcIhkk7Zh6ANGUQDg
xKL4ybKNvHWVGttDp85vwE5X00L567VQVGgiP1t+Mh6N5cG2cLSMFQPxb8So2a63hczfj8ZskAHT
FXC3ccb3S4xawa0oxCIdVXwnEBhTa9cErc8K0uJhb0zquj/zeZtPG5Mq/KRpNFMXX4KTM8yTkLFE
LcVdBCAIj27BShwm4CN9IsGn1FAVRcykd1XqHwKQiiROTcIpqmk57iG5wdOWtiydw/YbG7ghW7aq
w+yn28sC387uOIb088+xaowoGU4ZtfO9mApnIfVRiG2wJuShOvD9Ijni1IgYCDFCPfnedWMYNQq2
PMMqjzdSUc+6OsgDFUI+qTrxg/r1xX7gVf++BfZlfp225rY/se5F+OFRP17pmN3fM7FqhRRe+KCv
Sobve8zLCvRbs6PmRjAEdagDq1yODRCJFQDGB6AXbLtT4lBYyvZJGuyZP723+C75GQB7ZMrF1fi+
gLSmrfun3LVxHszS4muR67pgSqOYy0ubl1Xmi1H1TK+67WhsYu+lAxTWStuk5pq6g8D3ivbpXChV
P6Sy6SSi+KB3u8YskiBvWG7s1YG4jnfstWCaKCK8EJmLnbSKbYl2CCep/4kNCvzihdASCOB+GYF2
PVVqTqhLS++8uIyYvDnz84xMNRTFU6uEiZx7cJehvSe/DME5MBESptZSxnaLn/J51XDdOi7JH0hx
JC0Ht5F0sdt+MlYOga/M9DU5aGU/slUGSlEVjZnplTH9ktP/QF1pvQwCQJcz75aH6gHuM3CN3Wec
BKlOkAFg+X382Bjd98x+6+OiflLo0g3q2xycZw1in/6HKwRRnP4B/xcHe9HjtFwAziAPMgfqWqsd
a+Hf8sd3VkUFl6LVRhIlOZULfWKX7BREji4KN99hdGFSRDn2H1n7O8jWkpnGr79hAcXOP9OkVc4e
cdjWGQ3jzi4zs/bBgp173ZZRID9fUBZFXKvHzV5ss1nFXxTxceahTv/uW1kps2ldebM+c+9rm9DJ
xgh09DSFiEfAR9jFggISvX5lCQOUPaSabKhG5SN9bYJpbLNi/28ZQ/GCiWWO2eUSN2dEt5PFRD1e
M60F5i11yS5kkfuzHecHL6wNm0mg8slqTyyU/JLTqI6wcf0lP43KSOczE1F2vdWOW+I8gyLNm85K
BOhGaPAxDEiQPbXJ+FFYqRh2lWPWlo+UQ3WEv9N64O7vebiRvdWx+e+0rP90p72+cW0+ZZ43VC+R
kAeSx9Zkq3lVO4KusbD8bEQke9xq7/opuP9PZMm+qgYKKDTHWMJv94exK9PHYwrclILMocy/f/tw
h0Pnw5W1gjAMXffD1957pA2ZJF1CFMlDG/0Da3mRgLodse1TUQ66H4kMNhjNVwo8HiAqdA51MFz1
3Q0jnagofJSfiAoEKwh6VJ7rffZ3bDpjlZiB0PvyN4XmtbsGJ/M/Uck5DUMldZzOMxf+Kprp6WCN
Sg1YLbrq8Lri5FRj6gEYcKE4LIumjX+G6qmPEPpQZfYZzd26Ha/+EZTWz8unWaWdTrMlo5/HaAOh
MHRz50hjdQmR1V+ozNUy9OxynJSkmvpcKlJIGW7h2HVFeTH/Kz6XinlHCGPM5PxhmXZjrzCGtrIh
MDI33AKxNJhVfQXPwf4eFERDskMU382+Ea0RFQix3qipWMbplesfGG2FVqiEB01t2mXw4g2+FNA4
jbgY/rbu/h2dffc8fyteM1k3wItWv6P2FYf9Vjd4hdGxrJY3NPcQ7dOe8MsCDS1VOZO2uROwdrY4
ogRuFuK+/lZ4XkAWzd92LZNX69+pXNPTy4ef8ZgioRXFsdnOmSFX/w9Ai1iyhT8KB6hF5U1rCVgW
wWChYzdrMIa0301spZTMJxg05XVj65w8oAJ4TR1KsAZ2qlpAgW6eExoe1yAGsZ9xV96iZxvVCD4X
HMP6uPVtw6tkGFkdr0qQ/RcQ9WQACe1WLLj+JSOBz4kwFqBveJb9P8Uv0QY65CRBZp/nncaDcgpK
mLRY6enFznA7l1rmnDddzXzFS4UDsq8I/Hq6OqUzVq/LDdfqkwGTAEiHIaD1GRD+rLuzBVBc5kfD
Z4rutCi6CVVvbup4VGVIBWEAalX7QrAAwedRqiPCofLZAp+mp9rt9T7SyPFmM4Z1/KkWD+Tdyj/N
qVkZMF3balP64runLso2u5wGMAVFjiRpmqJ4JoNXhkElNp9SQFCP5XR3mDlxXIXcDwLO8yZZy8nu
PAi1i/nfa28RkH12BPUdbjo/gr4PYFlICUlFD8bHaL8d6X3H0DxrwtSvun6jm/Kpltohr0wNMS0Y
+0BJNwBpHuMlnGAm7OsBlogkUbG1aq7yfSyrQmotVglmnp3zunuS9VuRNJU14m+u/uxjgN2SGydd
fjeZbiS8cd2bwM06AoscaedEhFrxaAihKV1Bcozn94UwoIrm3mQygJu1tQeYVzZvFfDF3Kb/2TBO
3nhCbzT+xv0PRkYT9UcnxCRzdy+F/O1QG9pJYu04ZdOMq3/fScwiyl/mvJJn6mfagiiMIkqYrcn/
tv2ewf5vz94j4m04o/C9h0FG2VtXwX/JzKZXXOXK18J9iluuVgBHonkGSrN2bv1bM3kv+6VQ6cep
LjONTQxJwcSQzW+ISk/V4wp5+1zj/ro8iGK96R/nSnBTsLd+FpLO1cW8Qxmoi4cEAHE+AhbuxTcK
WP07uK0bctHIxfnZDXJSnECBypYevA0uSjQaDYWhJ6maCXD2IchokMbPpFQwlb5kiyZ7KeXqESx+
rFfNq4b0mds/v3KRKwRRQWJYneVLVJMwBxTwx1Lplvz9t8Yjk1IfT8101guwk5TanbP/QAsbLepb
WPO3aW6ZgIcescaWhAR317R53ooXR7t4zU/Ed7vUJL14fcHutqXZy8yIZIRAS3P4TI0m5dEZbdym
PSna5hyA0Xrlqt0Z2dY+eUVz3BDgE/e3Jss/C/EO5rQIhTBPXXNsicgWVHdimMyG2IcX63y5f4Ev
bYClYz3U86NjkbNR3J2Wg7mRHXk/V034ckM3Fsi0bDXLFuZXQjOmWV3dDpxB8Vfw/sJAw6z0IzG+
MFQdv7nwq6OvGZTZNfouO82uGJcPz4+UEW9r7qrTcURbvQvYMl675UrwFDP6OKuIYtomvC8xxFkN
weLPfrFmdoFxHGMIn4sZwOR9A8C11PEBrUEZW8oWq95WP60yQjtERnc78tZ4jAaM6jh1S4Xl5srN
Kxh7AJnbzPx+i8v8rbVe4X0EGuR5jp/qVRUkDTZd+fraVd1fhfIKNB1eoSprJM3dvhmEJfyqVtk9
rBY67mgTjW7vpbC/Zvqq+uqELPY7XLCqRM5AtZcI8M/i5LVQNGowylDWMWa0xN73jnUwduIRGdNo
9I6U+12x9M6JJqbwH6PJTnI2+vF2qBDWFVZ6VY2XlVAK7FkgmeULcGx5tItcbtFRjdbshRMFJxvv
DT1YY/Mee56Ido1GEr7Yc85lkJVOgt27KyYIhrDiHX8D324UUEYTfVu1kF4KE7g7HAPf7KAWbVp4
fqvOd3RXCWrvLkkucXx1KQT3y6ay6hBlATLoP3fnjicImcv4+58xJ0/0wDoco1x+EbodxU3UmIFi
jamSiPI5OhoMevYE/k9Wm8aD98mm4NAv9C6Bb/7aLOofwMF24M66GICdmeD+0Kei89fr+4DISbZz
sBtK9sQgksZjbY3wtE3B74r4N0HcpP5j/Mlff7ycdwfUdX478Q6wV/d6U8CKTlpIG2o351KWpsUq
2aUu/0u9x2YCWyct6YAYXutR1ixuBtAquJNIj7h3hjbCwejAtsxfoMEfykNYrC06aP5hrD2V0iAk
WppCU10LZSVAqQtrOMXD5Y3SQvREM/fJrSzU+chZIaYDw1ASglHCtKWc6syjASY195CDQ5vY+1zp
TD8ELwP+KQzR9WGnjYOkCDF84IHJKU6aeMQ1hGbpUKs9eNeD0HjprYkyRDnyPgQMUmpGK/RVHpKF
wZhpq+h9suXuzSiO8vkKzxYIueJLA/9q/5x1Frdde7qRL1ETlD1jljKiHIEhsQcjln7UKbyBEQ6O
XAceypltS1fIHSyx7IvxAsonzztNJ/GSYZuvGSIyfTZ4jXjYWTR+XPk2hc1UGX6vbfIgxtj2qAwd
Yh8zHzvqfN3hScuQ4/njCJAKYgR4z3+CG0RpaAxt8H7MFp2qTAoIGIa1TRzGsxLIv3az8BPlwjga
PwELSlf/OAc5CbXllbVxHqZvmuBtRHx0Wa26GH+EhBDQaxL91+rGG1DsMNDO6/0lbn5kAHvRmnCq
0JvdwdvP/XIRt+UfsnLHWMIiZ8JfPsR2+H9L0wiQBrYIVlk/1e3vF6uJIxLm/AK+TBUE5nWoMYIF
rN1T4VuXmwQp62oq19eUlSxOEnKCc2sYZz/ClRASK+xoG10kre1KA94WiR3ooAwZ59quIIe+wcs0
Akx6HypjFTlOrNN1qK0jP9FftsA6k9cmzKH5J+PRWysSCbF7dUHwhyxxk2ElW1q7fdQOipUfCfzh
F9+6d3/YFWn9KPeMSLmBwdIAwwxQTwKL306jB3MHj5LwJcqOTr0xYbSuPsXD7lxhqzHOxigtkVaD
Nku63fywoakfqor/peG4PxV82Hiqr8VG9ezrbViXziEor+9JbCyPxQ25waE4Fnv4aTw3HM8Sh5d/
SnACF5IkR9gpj/qYwt1ylasZiKXKJOp2t3zdLRXZiXIPSAEwDpshQnk2Zwc+Jgtr3mpVxY/zqwY9
LxNrfanYKr85SlritK0yMkDPH+ozb07IYOjSvRcnQtGhHkMSSuCv2wJH0Er5t5SVaAnPnYK7aR8n
InaAHSuOOcHSHSHn3FOuUAwJ5wF2fXaHt5LqAuaBu2C7QU8865V61DCq0kQf0kwtefbOwomj8WIc
auqBZSLO52vg2PPULrn5ebewmHaWxZZ1gBQorFYVF1mQGG8KMSjv6tNzy3BfaURC0874ckEYSDFD
a79r5v3yY5KUItCnbDTw8QQq0L2sjuL6rY4WUdgPPmLKcxE+vpcqVfm5MP5zReDda12gTTmYESB6
8LelUSwQeQ3c9XAviNCTJEJqcsdLa0K+3PrmyzLl93xMNFn+5iRT/nImSCttvt5CQXcPQf6lt/4j
1gMK87ZhVUArJ6IRxJizZWZZ6iLgeTtWy9KsbOruq736/XIqvGB9Cn1ZqcuUl4Ycnngl/CCt2iO6
MpuAfeU5yXXq8Ya7i11dDNpGQKH7zFEaPbaRCbix5rXgDEVry2uWh0mB3oGdgC3LhLgXZOSJL4fH
Xb4+RdgWuHApMdN2dRXh09u1REs7H9XwJrczc0/+yHpps1HQpypHgWlUNfyvtTbJbpPbAs1udHnG
MkmZojX6Me70XP68tvfQ3V/yXBWGwkoJ6BLQ4c3sRlGoAzFibFcPO1/KQ9bbAmmciABzq8aed4K9
qXVt61WAt3qxYmEdSNOjO4CwP8w1Fd03DfZDg5eOPfWLuRoBb0YyORcxtDQwqLDPWdPgUnIUonT2
4MfmphHEZYRfY0HQTWZv1dAkn6jMrAocyzT2e1ArhZ56UUqgZQR6fXaaKyY26WQCijqs0xUsrKTk
D0iQ1Om3trHUtUjsx/auSLPqbAOAH6N1ufi3F6ON7pWKVeD4yVrGhhS1h0b1xxR6lehNboRtAD+k
UiA+2EDmh6j6UQQN5UbJfdET9UTl0qusvXBsQ9ioemr4QyiKrJtyZzSinYE4PXKIotbm1lGy/myb
ysePrn/8A1vbzdIlmzFSplV01hUtuebrhWpOP6KjhAPtsD3/iDFOA75EnEp16tVlNUAiTpWL8pnc
JqA7pteawCUixmM8YbAaG9u8v24ne/jveZcQD0qJ+pfoQHXX2huIO2IeO+A/6eQWz52xUBNN2xdv
CZgfOmZ8iijB+dfwMlxBu0GzL5gMWnx/9dX9hKViW17sGWCO1Go/hwtpq9OMdzDiiAUjwH7YFnuo
+lP1iKJE+ltFRtfbrEU4I9MHf9ZYJEGeONs5q6y2u9K+eI1RRX92B1val8tApqklDX9ayrMA1TfD
9pTaXSIY67kjXPMUn3IxhMWvEC+ne0gTGbR64Ff3LDBXVSxiEyr7gL3KDVmMnOZVKvux05VAHyAn
/cbYz+D6lE5AiyRO7Vwo34Pv0ndAGv6cketSZBgOeJeriw64YPN0EcGa83SfEuFisyC1a7Rgd0TN
kgRuxJ0jrlLZvBOK9Skco8fJ78LJ3W6ixfZmKVhCgpSex8exMKCCiht1+o9WG1/cbhUQFLxVHwy6
hdY/1NV3Fpy9MW92x3IYvWkCD3fU1LG5Rxg1ZL/lYu1W3GgwmDWmrqm0Fip5rGDGq2RJBRO5Gckz
6ifGQbYTI50/Q6oRSj4bJtmRpG+jb3U5jDk31uKrpsVRXmlgfX06aIZ9fQDO7/MnY8M6fgpvF7ur
9iiQKo/jdSd266tUEwg+h49G+XfkJeYaZIu3MYrbUoAv6mSkYeTSPu8y4xjPJteHyi872WjaYJbM
H3ZV0eWNUBpFX5ksPwRhua+mQY9P1qkCAprNQ+EX5tqZ+V6XwTbGsz5iPo47jiSBIlhLG5UXl6h/
iRtU4aOB9IAX54OrENLkoXhFoLOBA4KUaIp3XT8XvqY1FSd87A6jPxyjtt7to8OdwLwDAq/+xH+k
Z+xV968EYxaBiH5vK3cyMfETr5GjC6RM9kz82Ranfj04lRposRKVMU+qVWe33d/6eTCm/pEHrHI0
kvhQopER/utnXdUCv1qkK0mrtwzoVFy8FA9nK6FZY4bf2oULPfs7piNMB9EOmu7PIi2lw+Dl6khY
MoXyL5nwbLgvU9J+0oVr3lg5bNn7I0kxsNFNLoFa2ZygEaxXICyUXWW2m6d2SJAeRte+UOGvft2Q
ZuttdpLK0dAVC783fmtALjzj/tJCuv/vAQBsSQGt+VfTp94SGpRIGmBjD9HAi7p1yQv39HsjAdJ2
noVHwv/ptIoskhzdLrW9cUcu0OgJDczc1EoYGz89VSA/83d+wk4WbT4+NmEc2lEfRSqz8JMBmlTS
8g4c6EBdRLsjsutEC/xiRIbbvWPQp0nkg7qPuCv0Zh2MmU+xcd6GuZirwe6G99EuGQc8MJLkv5P6
hsROYYqwTIXE9c4vYOcGRknJoq55naLczYNWtH/rS/4yrnzsJqhQTv4xy8fIU+2y63wPjvq7dEaK
zPl2P3VA13VRsrgcSWfPnhjH12/Cgajqdd/SurIIJXAdM36t8hfNtfwD3o25wIvyG/L5pUkoCK8/
yznzKHxrn+uaqrt/89iwVNG1ZKTjunuAndu2qmWuddecvERMeZXvzChOQHeUZCn9vEbTkxGlkAwo
pS12bDWICfP9KSJkayTGzL41WOjeClbORj614+IOkB+yKIyHS9VmaHYTj6kYj7a6WmUZ145F5gpC
bg7XJpi/FvIOnopTABmMq4xmApuSYfA6bQhM3RFpQqWrBxaU9P8uRzSkMDfb44yj0H7g7T+PyqV5
z3mnebxitGSdtD1ExwUfGQirSfsEtf7jpMcyh+tRwRDOzObl8qp/sEQWHR+xp1sCm7P1buP3Tnjo
G56hgw/IjZwXFx+B8Pf/g2W5CsT/WAO3S47l9sE7wyoRELFhViEcgB3Nzi2GcEB73FLVjCQKIAis
RvdvJxyGcKeWVWmCHxy5TapLtLyC5kIJFEWyHoNx2T5zlw7J+o2Ya7DFEIYqTX2gVAz7VzMnVFYr
8PX8RVX33TSqLxUtLfYhvRKRAuN89koFV6KF/CGTjIBdWjKtH3r6qvXSJ7kqTVKjV9H9fFTkW19l
A94HkrfGzwMeD5NP8lAc/kk1Z71kB7uUtWG3gK6Zv9Wom2AmINjivWEoIvkH5Vcu4uUTCUCBeo/m
7vAV+EfUvbfexlonTvqqQZZ11CZJtRICPDG7oVxCLrxsyqEbCX2AStSK7sfV7JyVT2Pxttaho4Z8
CMiOIzXfIfpEaXhfc636xsk+IkACr07WA9wI3mH2S49cTthwjGAfZeIjdwOBJyIsCggh1HgRf3yf
8PanJ+6wYMdSc1aaXu7lUELMpVr4gKjPai/cTxc5AAVFz8QmIy18jq5ZDCRB3dy+z3Mm7bMWBVEs
noMOdPVx3NNe8vMjcYGUORiVV3id3fCtBJMOqd+zErOlL1N0dnwMlRnVCZjr7VFmGyFNSEdW47e8
bDnMijbQDzvhDGGTElLqorxBkWzP1Avrbnt/12rq0ieEdwVflUACrsePVUHCAzDj7l2ekCokkD5I
j+dDTGLp4pOIiZxuq2WqiBatiXI0wVZ0NIEu+9gYbnrOdimAFhF6k2eJcJwqlYcuayMa6M8WaSFg
XyHgn4WUbYlwwWVA2SFnmODcSdnCwSHX1mapzfxLLr6xw82ThMx9WSTOE/ieeGfn1xbfIUk4qDqr
f/5afiLa51cdj5wMWG316NKX5WzKgn0VFHtOZJMTzcyXNG9I3w7vBUt28kpIgxF+qTSTn12Q578a
TpmNrv4OZtVmKuJrwPzHIQXvUiJZaEcN0BqDl56C8Z9vKzsR8AefbQrYZQcJFr6rm1xYZMvweYYI
vVxQTCXJ8U8CNBH1Zr7kBFpUkPyqy3c6HOSEbLM+CTUxRCjM7Y9CbIQnI9w+DdTSsMfMLn2UGTLM
glOa4MqUB3CFBoZVOUiR7+eXroYU+UB05Y4yTM95z+OmMzLvq3MN3r+snfgjpi7bEOyCqxah/6H7
40KSKIByqTtugHu1GYGEnZXsnUDmOux6LLMH0vmuJ9QaVvVSVH4tt24N4aCBkGutllrm3G/F4ts1
jglIdz4wMBKyXpQo/Xl8ZSYSL+8oCnfwI+GSVac0fEH2wk1BIJIAQVEDkpZ/EokboTX9a9GH4n5I
7UbNSFM3hZnvkTl5dIgeKdh0ptbMlInuhtA622Si+gsjpnm0MiPExje1/vVcqZa9bB0A+GUaUdRa
lwZxR/jSmlWTFqACSOJ8EpqoxfXwa92s19R2H6hy/P6QwrPcR1iN/qRnInltwGIvH9CqRnQayh0R
V1dTeEtgxQy593I3WSEiAmECHiVhmBGTMrsF2KTPg7zwgiyK6B+YBYtLyvxsiwXwbd0cZQXL3lXg
iLCl8DlYcKBgXvdq6bzH9gPIBUC/E+jqzITP5ZZ9yoLiXhJaVWtQeXpjPgRWtwSan2bnUGrgL+rV
URIjACw7X0rumxo7Y02C84v8lf21OSyQ6mOSBSd7rviGu/Q2VX4tubCLoJMRtWDPJXnFVMbnRux1
zlLdOx63pJ1FIwZoD4lqzvF9fazbCd9kxKNAwW3t4SsXVbfnjGwXPwnNgVZ+3c5US39REDEt2Umk
Uz0kVZ6h7BWCxKTr5Uhv0JmgMkCF6LRT4EeI77m71xBTujAKROqbvc7uTD2yeppCuw3w9s0EznUy
l3HUJoY60qFBa3LODgkZzTBcoM/LKuz2z9zReiXGgZL9chHodaBdPXCHwALZMfYayp/hCL8ahRKp
SzyepeeVyLJaGRWrFxHRorS9vhEWj85pr/t3bixfioTWuuU+JIXN2qPPFzGCgSDTrqk8S/GA0QcX
TAPF9jZYyr7kKjFZ3Yd3IU4tKme8nS0aDnhhdKWk/UnTWVWDEO9FsltvE2aGVgNurio740sZPryn
omToCFfi35YzYcEK83gX+CLli0RW0WFp6f20OZvB4rfbEQrRogUNG/s0EP1OmZg0uFkU2imsOSKG
42sKefsL/7fILRm3RnOdt2nPg7m2yUFm0dvdjeIzpQ7WLdwx8bApP63GSgmO84rwfRsfcLTP3O1F
J2+Nii855ltC3jf5U4bwy6EdXkUXsW/BBR4wzZ2v4ha/iQ7+EErqAlZpoQtgZ5RqClYysSuk5Z05
WH3vSr+DjWFsxxcIkX9BaOIQMuzK405T/MM/Rfy4ApDCJlQLR8OQMJnAihwOzzhdKVbskIaaVV2Z
JbT0K2N71VunHgWoaLhgX66WK/D15XJbp6T1D8q9dZ7aB7OIKUvRjW4ELY8fhdFNk8gmUY3QjVbt
JbN5B6IFR10/9BmyjjSM2hcwFIe+WxZPyOq7PO9976Y2ZimEwgdDTG3O95q8XGuVTyRYGkd/833Y
XJOg7WNEPwNdx5gw8Bbo3Ow00Z7V5tSGhjHvwYKnOjOFZ/zisUqAk/vMYIM7ixBfBkDKs9qgIm33
grOROcMobMTwspl038NU4vWO2csgZoT47L5LuyZEkjYEc2TBJ3kMNojs5FFH7U20LLDUtecSz9K4
GLyhd6Mz2RDczwF7053mVynucWrf+lap0UApxoDviLAfyaUIHVg2kiZYh/u9XPC0W0NYtNNosUNx
vNNPIyve6p8PuuLHa8hD/Uve8EA/ADK9Isx0D1gqCVd3dTcWuScWQBhpxQFFYJV5A/UxiqNcdmOw
sbG1Z57mrjw8dD4aIA0iDxE9Pl3wTYqQxXftIUKFQ7gexEQrtb32a4oTz4SZMFyinnWZ+KAMtnkL
9inV/x9ExGNPVWA74DLdB8DzTV/zC/Sqin7AtUG3TqX7v9YicwuBJrRAt1cWWciJLFYRmmAYAZNn
Ta3qzTnjvE8ElQlpj8Y+kMkBz6M0aKJC/2axQxo5BrG9h5O+nWp011wLT6omDcKWKStvGVIl8r5M
ponb+g6gdCAu46MW6L58e8GT2KN1ydSy8KiVt7DLKdUpUFL80ldaK73uPag1Rf17hLrXyEvAAKC7
knAyPNyCIPLYeEVj/XIVIrSNLvhYU0WNAvLBMjb9DjwjmMPi4WYJetr3J9BqKXDdmRrs0mrIg3OD
kpU0aEDzJqhhMLfZSNLyhiOUfjlshXlNxbNxr552Ep7HDErwFkdfB9Ctid23SQisUnYu32aw4QFg
DvUMkUjisJxWdfktEJPCshqivytkKa+iYztsd80wvfy0d12bTouNYI6bUTSaC8G+OrCZG67X4fpC
Ksz95q9Qmn79cXXfd1iPT6MVxMqEgfmVuC2/qpPCZm7kKfniLYsFQz1Lzcy5ewCERsLvZIMWrzwF
62qdqfutkg68vP4MA7nRvi7bOC3329ELUldxpG5qALqEzq0rMIt4fAO3lagzk0Ks5MeZKB1ckJ5P
nERU99U625hjgVjQskfQX43o0urBiLkWAyDxPCCBhoZ3ZSjmVuJ04L2AhBZGxVrVgTn34qNReuR+
pHhpehlFJZpUcCSUeyffriab8KeIvX/COH5daxYRrlUtFn9gfRFgVufI8c792QUU3VoqLNpqbejN
6Zob7+R0JrJX1BNEOJI3K8pPMKbkAzEaubKpVa7RsrqXoBs6p6ysdWhGeCVUUKv+ZCL3+PuS4SMo
BKxiA5wkWqO/5B9AjbgeivQVpzJiOUrWcxK3810xFw2BqH1/wMlMwrJjJFINSnx2gCKL5Sux4xxg
L8TOwNg/LxQ57naiJIzwD3zki4FXK/spsVr7O6sNjTy4YSwR/VpNmOARss2RwPoEQy57IgcVxIOA
9REWic3RW92s0scWCKzzaPWhL87Gt6/4KBdVYSPTq9yVcIPM5144Xwl00NXQ58RYWFP1WnxfNTJD
yklFMd2I088I3kJ3aTwYdBs+34SsUkH/uSReuYbFglMwL9ce7qA112LDZX1VowjsuBKTni2YuRPD
zC6nG0Iwq9w3SvZ9uaUYTPz/S1mT7I2VsEahYcrRuvbmoA1zeZXWvSKs2ZEvg8xWL75lMNDF1kzg
ivA85jf5IBLGreqywzzjPVpxxmBjWK01IyFI4O/3pt0rlE3xHtArWgp9WqpNsO/87A4xObgi8RhD
ChuIndjrggbOjUL4KUEybnR24X+kC/yDXBOB1A3RefivxOzD7eFvkFd/m5FCWo5HWMwzaweEgWk8
Gx6AqJv5tU2BjbthL5feV7WC2jJulZ3QazFJTLBxpnCK88LI/h/4wjhax7YaKioFKTO8wwZreWyn
RWRO/wwLpq+nUd6z7V8yNvXevLiwX9Br0X3i6SawL46FqF3cEEtUg5fmhHAfmXzg/D526P6HpSmt
384+Fe4AsYRKeTiq1laq7MAfUy25mkFk53FT6BODzSUsanHeaZmTR4DyPGvJXIrHket6hrAIXcu1
ng8hZngIOqBoD6vfwvyJ/NYJj38v7Jsm5Qq7Cn+MWQdoHIOE4JGoqBlI6pb3CTU2G8zOFI9Xz2qv
n1W7jw+rQ8S2xxt1uByOBFsWljCOqI1T8qu+MgMW8eRR+kIY6ph0cyvXJm2i2A8AYHPCKCKQWvYD
22NhKydYZqT5KsQoR54XL8xSFIFTrWjIDMRPiI+jUsMsRqbYBMS7ebVAyQc5w0dBMH5ULa4N5Mo+
ziKQOSaeuOacvbvqVRAnsWPraMFn7jMJAXsv6/mysHxJqyHNDb+7mZ35MA2CX6TNWJnSAWRGvcvU
YIPePWExhVL3D4YT6AAveC1vqNQUMMMDKjgtLVzsEYoffy7loYVi66+JKgPA9bTXaP2mk7qomFVr
tOL6f6F45q8zOa2ErQdsw3MLk3n3/c4R8ek2buCSGdZR0t5+PFfDoTAeTqeAPBsN81l/LkzfPi3D
0Do2IZq2LTsuKq8mKx5pJx9HPOU80B9bprDepNBit7+52wu2mOVklojq2Vx6vTO1WIsQ5R0+O1OJ
9Ibvb7WRYvoK5BI16ESH3mslssoWkyjW+a74NSWvktlDVN10ylPzjl2s50RITmO62dNY0QNoICkR
+aoM1fjWaUIzmh6H6EDKaFYajBGOMaTUJy+6F+zZZL5HIfiVQFk3iLR6JTUV6/SmHFsZ4YoBioYx
Fv2O4KPPCtO5TgU1+6vnxDh8n6FB98GioG1Nv/lt53tA/J+p8/UxG/EUWyQbE+bUzMOqtHxKKhvm
VztHQzre6aktgRTwR1fi/2udYQHCVwfyqi2Rq5T3KDEL/GDqK7id3QWb63dDu7OLjof0CcRICMlF
ZgHSb/HXIDyZ4McwTjAWBjmblkThvXju2RGesMVmLl2eEOtsgOU/U0OL1vv1y/8KHljF+9p8nlqK
0rXMs9YjQYgw5quCWyiN9XZZnv8iyuxQ+Tn2KXnz0YSzEYoruL9TSVBtbD6u4PwXe73MuBIKoiBx
4zKKSze7Gj0Wh0IPnO+QDQJuMeQjRqPlmOkOuRJADGhjn/isitFSWDJZHRdHTZqP7T/l4lU1WJ3C
q4oIxtKlmhJLs6UleS7onB+IBKBBm6vwmMxH1k9NGYrNslKEnOmopSfMHjwRTB0EOyoFETMJDKAo
/ZrYUk7Z9i4Z9R+5MFyiaJ3OVjcj6HyCq0MOveCEu+o+9Z+7/YxkxbLceBVd+qgwnFL6iluYZJru
tSjXL63EKvoUvK4Bwn5EloKJ36e0Z1Z01CYXmBfPVbGlrhOk6mE4x0A7MoDaCkJ238ipcdidBhn1
r4BvYx1pR35ccv62O5W5zIqgtgoEvJbeMYguA1DpwNK0Hnjam7nD63+B03TjnjshgDS/H4seJbXh
c//x1DLNa3wyaF/IW88V9V9Skp/GKASOW1H2BMTt3XX6TwOTK0+aC+Ks4iw4j6xDMYhDv8srZbhP
fGvM/avqeXpj6dqbwV4P4XYjGaOersM24PbrDKiMhcpszhb/slZM3nEWoEENh7pmjaTzwD8BQAlH
ogSophXsCAPyYQZqYF9WsCf5twLDtq2H2K0BgoMGMjOixsmHUfJ62RdyZisavHcCTSmLiX7bBt7+
y5e6xnv11el6V1DiKQxYxUSkK5pssfVm+ZB0leWH+yb7Z2M3f58CCfCQpyozmWDJ/Yp207YF/WPe
HOyuvhjuqc/wAddha9/sECKetvRyWI+VYP5H9N9Y5cqQ6pki+0gccRyFOvzlRhDgcMSQZwW6ULm7
eomeppaFqBYcuS3ZA0A4PsHfUl2n8UGExbq8m1wF135dQ8Dh2KDQO1FFKJ5QQU7lF4uiaDOzbtEF
QlOhT7ynrtWGABp0BYv6giSaArOx8HaBV3a7aw7jXFdJ4rjKCNK8VkoczBd2jxWtZE0adchWZ/Ud
/WAQEIh8bhCj/k/g5tPCqEKCJao0vN1yy3qGkA79YjF/O5TBQqcmimRHZAJLAzXznYx2Sz+l3490
v1rX1bymgscSMZn0DM8QGb/n2hl52YkbAZd73hTNgwB7/edxvb/jbGledUIuNobH/Y4GsinWnyiN
32qDowsSlKJ62Zusg3+fyDXnXWdAV3r1uw+ms0VKq6Byz2qn3A2yPTryGTZvZbLvRgMvOg6Z2tFT
3mHrWuh0OtGPbV9Imgz/Y4391Xy7CgecotrEZre9RXOnOLzn5iFFFEmFyCqje+JPX0oIOeN0Dpe5
/jVwomZLC67YGYk+v62WSq6Kh11nPb87cOgaVNV0cqMP12Z79qwkv/aYR7wKf7sj8NxP2lqLvQrx
pAJMEoaOlRkiPsQV9EFUhzor0M+EiJb3WWh5f6p4Oe74XL3vB5q13pvljYqGveah6cUGwNri4Bbh
5L2mXseLUHV9+2T6Qus+NwZ0mEWQWYelONCh+Si8xUjUA+88CPL7Qgxkot1FyRCvQSkohHWkaB8a
dR3FNhT/sfg/+6tpFo2nSre7+gMh7O3GiNB90tvgWVnqwz71RvC508REij1GFeddqmShPHslh4ok
lwNP1dO/xOaMlsTfzCrrF9f/VbeoI7oL2DdhVVvf49aE8vYwWxecY6ezqGwfCLi2e32PkCE/6MRM
hU7tm+Km4ozYJvdDUqQWzkVAE+i8TOz1idKspWT7LKYbPNEHt2vtjTLVsgpqNjfTkCso+3z0kDzT
zuxRR4yd849MMssrfDEywx8A+6DdIKi0xougZDzaapZ4bsKjrDfRXZ92EtAb+b/UV1D1TJsutytv
S7oYozv5bDpHRkDnqyN8B11hFrqbdp8ry8HXqAcuHL2f30pOtKqiN/mK95TH98xhnT/TLh8+UQMb
szgQsJdVzxRqTAq6sV5bMBV0iUILiadkPXQqN4a9ffwzARr8Ae+bxf+sBWivweQGiYdFkpuUKl0f
PZlGmjRDrvFwDeadrg11V7DvCUbGh76AgcWXMKA1H7acN99jaykCDQ5Cqgjg0RzBq9jPxFyMI+as
gqhgRHf4osCfqN/bGJUVX5KDCNhOEo9BNyZp0/n1tMcqgD9JhcdocOy63dpwIIfU5Rfmt6/1mdLD
rr7aN8BtRgjlJoaXB4Cug67kcLdyqEsyza0+ZeLC2b0TXCAuqJUae6DMQoa2+PFTdn8EviEbWxo+
8QBMXpBJISw865Z81AE6tmmqGptKP5RCW6KPbW1ATgLgyULM3Vbeevd93is/NExN3+m/o99G9L7K
R8dJQFBhNLDoNEY7egg9p9srvsbafCyD6rUTZvBVkCFl1ut82hpRDOoLu+/imbvFhkEp3k3ndYDG
EP7m1FXbVcF4o1aR9Ph/09s8Ys4i1hOYVBh2Q6Snke4BhOeBHfU5gJxlgPf8BkoBtleB7wVWsMNt
7cp4VdJJri9rQHZyg6XauOLPTGGE2Th2VWt2N95CXMpQsNtzTkOLxJBrW6+WlkWgAfkzomGhL3T5
yzhBODTF+Rb7abHIr4CNO7vWq45ry6QhSnhdvlIAuc/QLwl50rDQjLHiiyUWT47MKNze2/Rqs8Ps
gFHyjYvYTEgZWgLf0ZM2Grjp8lYEfexOy4ZK6Uj9RvKPJWc8S/wf+/aa6/HtIS2a4kQM59TH5OvS
hbdEVfUeBxql9uVlErqad+M8hRAkg52OIdklpUAAKSdQ7P3ND5u3zGUplSErVEY3x115Z57VOQUX
LFGatCq/0Iqrh/w2WXXcyVCZ/t4AHu494M3M5Ie362hg1WIDQsAvGX0q7pfs9pklNcXBDn+SZe4+
UpyQBPDauUUCdU1+P1WgB9CutoyfOlujRxLvqd2bFIm9fTeVPJ0AW1CSDiCeim8/IywtxiLD9MJs
r8yCPD6ZMM0xYwAHNh4/lW/LGXm70I5WTgZF0Zta5mbrihpe7C+XxdoxJmsd+8iEdd6Wr/693gWI
ynXTl+83BYc6Y3SXnIDkA/S6znD++F7rEc8Z992NWO88BXu42Lqx7jATkGZw1wepLT/mtvi8QJag
Lzk/RT0jsrOlubRg6UcR33wzj8kbOkR2nRo5ZJsh/yASy/VKtlyhU3+EhEYNNAD48RNL/rUPgdNb
zhJ+m+lwUB5W3b2+9nY8ECWgae3Amr7kNdKFcM7d7GxtoTuD/ddnOpAN+pJz0ux+BuSK/zn/6goY
33D3VwRBDynO17yf87J/LttpKdVQcMffg3Ey0nIcTkuSiOIZMfOZgGXOR91Igu4X5T/LhTGNcrmh
Gyr80hVLRCMupc1obs3UXBaq9AYcHUa58bdnHbwQ9LatZJi5sEdcDx0lvdwrlZO8vVA8pTLH8yj+
aGFvT7Sz0jMDGvGz9oT8TOYrdPbZ/yx47OxyeQfDsVzgFIfqzBpAEBUe4ZrEPBG7ixL0Ht6m6NGs
18wG9HdR05pPfHR4GIc3IgwzDhusQXcgpomRkOYaiuoTEUZGecu9qtckW7Z4Vf+p85j3H6F+gDzj
YpEOPmEdedE2xgRa1W3NrHDrwRTiaAXBLasGZt6XoXAwBpK+Br5L9CRv+rWOdJ3p41SEMAF1ZVqK
f3gTEtBqI4nKBdb9MJHBwLbhghj5mW+WLBess9OHwgdGX753BM+IHebnAqvZRkibyrcn8kl9Mqzm
gd5NKv2RZ3Di2W7Z4uvv4R6FuzA9MMJYaUkEd5BqUr+49ijmt67VgYIofNkWbhbLSwzF726d0ExY
l5WSoBWe7PFlWZzL+s6Cdi0K3bciaDRm/rbYJvIf62XEH8QpgZR2PMhD0TrqvHJ+IXQpK3r636mQ
7d86lbB9YkqwtWOJQvRApiyTCWRaQ7y1sftiGNPguNcmOuMr5W2r8ZP4fPFdVA7BfFeQG26Rl1KI
5QMOnnKSAx20xRTwo0jiHPBPshXTJJundnNlq7NCH7IEQJCb13KDuG9gpVmCRQPC6Y4vtc8reA0S
PdhCYzpN0vRDfzR9jAlqWLvG18JE2NCotG7LSgOYFIi519u78XzWDKShhapKD+ifBNC4oq0k8p/2
6nFZx/bAJHZEWho33pk9E9m7vSQL0J14cMDrjSJh3wev9zgV/AERRiWPuiDB5beXb6ZCYW+3ATbL
WqJjp3Pxsf6dpK73y9erZ0U/eEspO8QPuOdQNbAyIQjkXWJAXcA0oPIxsMAvgRnGYNH8nxFX5VDK
J5Uq9jtotKEhTz/OlInq75uz8wS4BMwjwqMQkvDV7x1Z+4VNEx8cV5mMEy0ZaRAA+wmX/RAlTFfr
njTDPX6cFWtPULsPxbxc0zXrD3uEcZRBXlk/CDJrRZFaoVqeJkCfInCrywZjnTXon4g7OA2PmiNx
9a39vbHek/71BmkkyWxsN3cOJUzQoVpfAu+wqy0KR/KzCicdQ8PWOrT4AbNr7S+5L9KZJVTQtiYn
KnhgT/Exbbn0WF/P9JGmruP7MiUoyMd4AA5FnuhNEvmlGKtGLepiNbqxhZyk/K6dwsBTYCp24OQH
u4VBz4K+1c6PnkXF05e8mFfBFqWQep/rE9VBm8BOBjGO/cfuxoKNB1VPRpbtUZxeZ6DkSZFMB4hT
WjtucMA9wqqIAsNvKIxZJzOj75IPEdCdP9/hsvQhQ+cM5hV5rP9Lb+P9UOsFaDgzaBwYmzmol4Rs
oIJ1bIbtU/xmMu5rXVCuB/UtYoZvjMJxPFh/Bs5uggfnnR15KylPEg/yLzkfJ8IPdQBHaUQtiERK
g/MMRxxTAyyahE+KiLGugC+5YuPRN09nylUYj+LYpKMnePP9r+xHcEtA0hqtx/ixPrrrnO6xIHqI
Et43apQLSjZH3d4HzCs/whXa0s806uPr+XHYO8NXN18ng+zHBftMDmAXYV8RbvEjG9YThnSd6E2h
SWN4HceQPhq7X4xt6vxNi21K+s+MTfhb9R1zqXQcYrBU9NGICxydqrbuKWenCOym2h7WMEKiGT14
0Nqx9tJ2ZBEoYBRs8fw+9ayZC18Kb7Xv7Pn5rWQTrnJ0/mWqK7epZEuy+SQ3fzYUj8IxeMKo33pt
A/FkIcp5pxNOtg1kmyHhSKxFBhf7rQfwAoPD//7RhHqAMFWMlHtR+DRlHy5MT97GyodfcTuJTkt3
4B+pM3kmpAxjoiSaS75KGQrTqgkX0n5AOzRY3yv+1MlYepgxRnbp+5GJN99Lb4wZ6Lkc0qtny5IZ
mfMImoKEO1XIxqd0opOiynNMfXYvTFVFjKSSEUC48B7yMf9N+a8rAuvKxK5e5dJY6l6PuDm40eJ3
07al5spiiWWyubOeRNSN+iilJaBmxcs+MMCrCFiYPpm5dqVMfpqXTVcYZHEbj0bLRjzEiK29ducs
yv0fp9Fjd0yb56DSjyyBLNA3FvAP0Grj2MnsQXLPdIY/nDTtTKtNDTw0qtPoxydDvEuvBc3htVnA
ksRZPjMJI61X9/BHrjvOP6PzFNc4uA9TwYJAJyI5zpfxVhDkEWWay5AUb0RqWuhTSB27PX1PFuEl
Rc3IDqQLtkVc9CCTrCLooHP8Ul+v1iSAopveNmgX1bg00PVwfreZddcyKuWiWtWQ05Le9ptHDUf7
hMY33CsWIL//ofFlkP0LV7/6dpIx9PpKab2a5V8ASrKhXhJoDS6tl+ffrAacHbHPanplBydElNLq
2QUHeJitC3NO4fpFkoymcD6PT5RlvUpa6VdoM5rg80YgGaQwhta/v3GvZlWN1w/7GhXXXAvobwDX
VOMpDhFyw1/Hprj5REcGBfu3UROauebex/6mjoYrnd7cR517yHVhvr8dCnMKLGoMm3vjBCQQuiFr
N3XGQEspqupdOnfmUF3uh+k+eNvitrrrhq6yuTmsJmKw123B6x3Baz1VbMXAmpwdFt0o+8N79471
ot+eW8wp7d6zb/iK1H972BCNJGTkpYyeUnjp6vN5GYMz5eclT8Y/Iw1dnbyqZW64FBSOGelafCRf
6d8jrBjrh/vagP6QgzEZjv3/9GqD8FChVDIiABeqdEgmyrlaO2S7YPW+QTPArcK3wM4NgGXQ7ITO
YPt4Fr7bJdfz+M4o96evgf8Wrtsl/at22uvJYyJnAkJfXeCf73im4RR8i7i/GpJOrERHA9uBaglK
oA++BVWeAC2A6vmsVDzxZrYON3xKrmw3mUdmPpEVRxkeSgJpse5/QEXE/JUaQXDwBHJizyY/9IHm
ZwLbb5xVqylI9XMl+7SZk1Ix3AWahrMasIHtu5OkQ6wAeQbSteQlmqEwvVq64yiN6N0l6wfGpiir
cs6ywpV/zxqkM5BfXbrgaeDOadIZxr3x5/HS/EEPaqfPxuIuC97W16Hahzs7L7iPkn2vDW30KBzk
D3EnUvoPyvWDqlXZx/7z+I3nPnSVKPwl0MFECW38RuGf+FNqkXmaUN3gZA2tAXLnO16hQwBJUzO2
+Dm8tkdlrI49aK+G+vYi6nUQKlYz0hIRfjw2LnpGU2zsCNbH+Mkr5jMynvDIyvWNjyV2i4zz9u09
A3nqGTljWNTJEj46iggQH37nOlhlbOJp9Qfr8JSEvMmgPiYGCVF9MtnOV9Zne0RvuYUiugc3T0oF
feyhV7Kxm9S0IOl5A3R2rScpLkvyaXpeu59twSHpYZ/2sL3/Dn1h8TX7tFWRUvnThvPxWFsWhQBE
8uOxj13XlWYoXeijPr/x6EkSTQWN2FfRalmLTeQJvaf1PVa1KgkPrpDX1qMR5cAdhSgOFPaYZOwM
RYWSI85FSidKuOmAu4m8oBC6eXySLc/i2Flso4UjPz3JMdgTwbxJsKdKPtsqKFzvr5VOQhhGO8/5
SdVL+FuNk0jZuOIOwC3MFuXMSo/FQVql4x3mOqc3+rIVDl93wIxouYCiHaQsVeOAlpP5lsCltZx0
GJ/eX5QXhxvvyFNTzZIXPHf0RowG54G25G0lDtu5FxUltzRcKPqfQm95yQmCQG47yLqQ0i2mD5sh
BhkEFLqx2zMoV9vBfr+OxGFTw07kM3PvcaJxRQyiFgj+cveEw8FY7zzcxEUhkBSwrshw/v9J1fhE
ax7DDi2N+W07OhVZ3BlYg+M/pVwmI+uroigO1zVWRcdBBDUvKj8eK03qyG7+/NycAluaEJViPj3C
ifx74xIj0ihEH5STbpHwD6AyxSWBLgQjsoFukqnVgM6ba4jtXoy4WNGwKbIwDrZowtcMgkCt8iUR
F2cp0prbHQcVMfvnK0+AtVR+WDg54Ho7fJkbnRNstHhQd0nrY4BJh1ZZaMxm0hcWghMNmt2QTNWA
DmL7GeFccehiLeOkeykh2/uf82EK7cqpCa3aOCFDztwpD6ZFL6hyiEwHcF2Fs8AEXUBcgB5q2zUk
Zg1+th1u2vfXwOUSEAzKtvamxzX4SOf8u75hGW+KHIVEncXDT4Q6IrX9/uXIxEjOwiS+eE90rKLS
GgkpKmCWXG4s0r6Sn7SLpv/LzWe6ZV0SkwMk2+3iC5BF3geBwIUwrfNSxH4ecgpMtuWqtJY6ZYB3
fF/MnrlfZUUSdHNv/wDDIySP6etju0Gezwqkk1DRqZoj1TEgbGTG0Sawso1Ljs5WNPrf3xOP3zl5
9512h92ZGJyURNe7j9/RJEZNLKJm7NurMQp9LhUWu7zZU3aCaYnxb8WHiZeOgkncXHjYGfNrFIH0
hMtkac5jSYb15VauVq5inl9qfxKlPrz62BSTJNVjL0qzRAqvzZE7o8pD2y+hsmha63xeSFFj/CKf
5LFMl3070WK6renVdVSD9symXYqxYx3xhTh24n4qIYseUsdwkG/Fv9njq2+OEkWnzx7rX7wFejGN
Ez1UGZM7vheADBfC1Thj8kN5OuEeN84iQxZUbbYJN0NAl37sv1pasSwI0UNin+YAOLlD5ShwBYwD
mhlXKf/0IpXboPdliEn5kv6stTNrez6SaqqkJ2U90FJnKyALZj+gu2p6CvxBWgGYSCdGvh3eLS5O
SFzLKcmGA2BW4rk0w0v455e4imz19aNzCsfvSfaX/jBuosHCWq/BCnUls2j1PVWzsd6bcZ8V99Io
FJpuHFUbsy57ibjF1c2yYU1eZU7J3ytsGK9XU4a9/tSoWWlB2FcAU4wkpmQwsLr9R9nbBmefQaSu
0UHgi1YUesL7twpBIXt4YQuBrsUUkBh9AAkN825mLpOWVpRbVEABIX01iOBNnv6XDmvOaG6Gwxr6
6oOhXq6ipQ+YZx/JdHLmxk46vg38vBljPDszzJn6tWn9GX+IcDyb3gJgH5kO8WrX9e9h8y1zCjs+
jX92GuwABe2/WsxZVa0g3cyJFor4XUXvlGlTWGXV7CX3J0a4dwsTZrssHo/tkQHMvJMuFzTjkGyt
UbQGLcCDGI9f6bkyCGLpo4658RGLsb07fPuYm7WYAucwFvqX4Kg+8Em39HJdpJX6mVLLB/catOeX
WbDwEa1pz/wSna+VH+MQl9VwpZgNa6dExjqdegdH+PQmZo9GkAa83iZr1OYpLNS3v70Jgmk+FvI2
jVko67T2yZOnPjhqhJTinnwzHqOoQRtwZ7NgyFyxikj7qHBgLP7lB+oZ8T25lENTHpQYu6P36myn
u4s4bnxJVc18C33R6lla8lP/p5liAc9SguEgjsTwa5qKWsNNSMeNmVzlTK617KvYu00RjbftA5aG
DVLH1L8zBrY/VHy5eH/QdHQFtIcMmNboK8TkTDY9+8tmMQ+ANkLg+zU3S+cxV5NQqWFNe3rmvu7O
kM5XnFZ55f/u0uEV1GmZevUqqRReEp5EsPku2ZmclPv9FuGh/EE8GQ4cC2PVooBbcMawjJvX+X5+
tBe06Bfx9XOwZfE1hfInEe9m39CzpnPHLeYLo5zY2l/gmXQDDMCVXt4byrOR3gztaFXsRM/F2Ya2
eZ1J9BV07tNJXpsh8vvlXMfxeMdF2KMhqFbJqluICaAbx/QxA1WzUUooX7RomOnyYwCxsWabMROA
iqFVFqs1uXu9fkekwoJmIPL67bobp9A+ZGFd4/oNAsemIpFzLlxPPsVvrZ8dSFu9P3B7ej3V4Esj
JR3/fxzwreWv70p2LpjFytT7bIe4DDUTXedMs65fWgnhn0FsBu0YPr3SHuqhC1/gLFt9ESJzF5Nc
TTMNLXkVgESbMAus5NhqvI+Oub5dSPDINNiy08hlFSTaTjvYeQvyk8+YUZdQTqoVw9iAKjy6ByZ2
FNP/0axaL7wHHLR64zidoFPM7d+2q37Hnv08kWS7qUgZM3Q1fetJy8UuxHiE1EjFXBDSF224tKRE
leu4L9k1T/RetBh7CrP2lhzPamj/H0SzdFq/jxvnJwPlJw6j8yQiXXOs2Rwy02GV/3IWBHlV5TSG
9kMpg3g/cfmzcTb/XSAivrtI+pneqxBEtDtC9h4rQOrXfAH8K4vRI3rpat14Lfaq9EXRLi23OBhM
jufRHbBFnUgBLnP8WdZIKPWDm+L49puOL+OlyeQDGsjanXHubqtC66kbM6lmj0QWJdcz9VNNaxVq
dtzugx9sa3FS7ZAMW0YasoM/MuixxapWWYvHFkQKOXohHJ4RGLb1sDIPLtz0Cy3uN4mjqxI9KsMb
tOHQzmaieijed+8T+e+T8rc+dx2wQoc0c6165Cvfk1+8VEZm2HoVYUoKEoQSUlFBZ786dprG5ldr
IU+IuLfbylyokVXEX1Pb9Y44LSnm9zJMxztkR4tVU0Vi2TQ/JcovnupQGvMnmdrgjm0riwzxrWRD
aXu5SavgpjbA6OjNGbuxFpzR0Y4JVhu2DAS1Q/xeCFD9KfvV9Z6j5pifRULM0iJE89WDx1wcES05
HtF/Iz4NzYnucwhZGVtmBPqd7fTDRg59KiJdSR3fxsYZsss/fNn+YkL3n2y9PQMvEq6h4iZTaPAW
fR5awdzGxe53K1NrovH7VXm2ePCwhW71M6s/s3qqwe2Y8z9E5B9ntgi2VqX+OMauezDnkNeHiOVM
7WHxZPsFFYN2TTjR31xWFIlISR7ifYoTuAcSzgG2nutoJR4ELy9kkwzaJf4ITHAdKNBJJlBgFsN6
6keHe4rU9VH7YghGtn18zX3xM9DWppDwdg15io0XnYqFgd/rcfeXAf5J+b41TCSKB1IIWGrEkTt+
EJuYlxCYlAfSxOk9+/WGO7n3R+kx6w1a51STRns0usraYkoU6xyatu76LsuNj9CG7kSJdtiLKvOs
Zy5jQdm7ijA3B0WSgVIXoRB4xlJ2+2qCWRYiY4yM4DJL2vUUNhewOtg/T/jQAYEdBpWxbEjqQBu+
JS3bTRV0UfMyvMCIRxlASSpQqEnJVeQdtnnMxmU/VeIekihOhUJvrNgEWjuqHWsvrEvp3HX42x6C
pYdGoUqXMel8rFq7nfa9xmlBnyPSUtYfKwwfW8lkE9X8Jiy/qQ3yNJDXr1SxEx3PXfikWVGe8kfM
dGI2W+DbQ6cPvh08DPgYchbPW8OgsaRjaCxR830pglGRN1Nz/PH6H2tnNiIv/MCuv7QnhYMhtVhC
gfQyakqx4IGWBagM39NV7OAP4y5iRtRbgpX146SjMCWxjgSw2s6RYQl5Pww2uUbzrCXgldUxiKrN
ixjWe0MGyBSlWY6To+Weq0UQLSDvnv97ley3MRBQqogIOXGqP2QiD3SFLMH2+JM6sR1+0sR3Zfju
wyk70fv4ysDQOYEKGNQvSkXJcUixsDtxdBkkQlPnqPXsIklBbxnC4uq056XMPBPn4IC3ImeGreqa
sJ+6l89ZcTx02w01r2A+zf7ngs5CH/JLJoeypERnGBmabs2kZlo6OdAWq/fCcG550/oLanRWM+Lh
dfN+BAHI1cXHzhlVxFNDdojNuS2dDqnrZ381cTp6k4CfiuqBzF9XSz7NrrbbUl8ulH/LHa/wNGTq
ebnxGWnLwVI/JvAcnau6IOq7Ve0TzsVRjCUQhke1loGh5DdcSN1TlvVImsRZ7t1HdBbM+9KCstJ4
Jp7+3SCyjqGVTBWBejizlunwoUpD/iPVe4LciNDnkCyQl8wotxO9XKLUllaQv9fwd7q3+vDqfuOm
6EPiLwb8ubecyHn+QwH8n3VqJ8xZsPoeOKmOi9xGsLNUjVARcl7avgEu9sPzJpAu4f9zHPYlhAEO
uooZtKG08T8sOuCSCdWMX1dRhOANFLYd8Qiknd1a/rY3kf1d6cN8gbFP04GnDl+SKUSd8ysm3W3r
wa1BXHR3iHrbAe41FaC6wvMAxhcVrtzTph9J21/oSNBPXz948hVTMpWfKJKE6ivsJg8ZdncCA1ic
U7PJ5onNMB0/7mFdvPNpXGbv+alhopgOB7urF7MyBaXAm+5zfoaemL0+DARe3fjUevo94Y0iDM/f
ZY2qUHu+WWh2NxrWL5RzUBebcndepJr58PSiUTK+miM0fSHqTdYM2T8UgPipzrF4orzxFccSaeaa
Hy/ZQAuXYKtGq0O5a5xDjXmUNmCDDW5mMHvl4xnSbDMbP1CpCMMzhVjwYvr+ZQmgsQ/PFy8nMumo
tvbC3SGyG3P2Getpu9yiKQnLOA1Yk0DOS9pTgcrmHwBPgSanDgfaXd3Au5rdtUvpO9zttxPgqLXV
zdf56Yl58t8iz5M9LkC5dccZnch5CkALbrJLBVRyrf8YZfHtM4ZbqU8X/8sUpSuxdYQD1yvByNNT
/l+9WuRpOdRygT1P0w+Jom7VaLBVYGId/usR614QZlzJvK2hcDqMIPeJHRxNJaVTIHvbDqV6K+IX
ziYLWimkMzq8jBkzyvwMDliW/M/CgR5ZKsji3x76zHHPSsPf/lbMq2b/ie8nOkJBM4gIbXA1hOix
5BvewLvfZT5T9Rwi2HtptnteRhiiVvCR5K6BnlSxUki63oGAn9ly6f01DJ1Akcg6eJCxD+8VKaM4
tPZRwuPk2mf19MzFxLeez0gRlxVbO1zTtXDESIBcLJL/cimgMpAUz53VKzYAwFRZdqUqCQgmmF8E
L0CypxOagY+NNJc26U3om0QaRB9f3TlbedJN/8VoHvq+bCeuVcnf485Yia0vps4SG1+LNcpQ/ME7
MW8JkMbYv5CRML8QpRuxLVLGPhuyvEAbAGbEyHybAn+j93Lg8QbZfDZTLny1C7JsKECT5Aea+PfF
/KUVxQg7/4j5TO5e5xG9lsMLF2/VhqJTwEk7DH7pgpotgLTICdWkZMmh1zewUT+6/eRkHidAasY9
jkBU8O4wzKvCTs8rchttZ3kIHf9TEKKYJuiaZ94X6IM0K4jvfj9kA37ODdFxWCmWvSnA73mVbgoO
Cw8KxCkhdZ+vRREpaUyRy87MwDvrUYEc+l+t2HR0XjorY8Tn84xjQacU0pB8blm+xvYhSriJhVlQ
4BUm3IE3ztMKpRdR521nhYrWDlpmfvZLGf0ei4hZMfRl5n8n6qVFsfAT5wW9evy9v0eSBrNgknMr
joxAvwaf4aQX3G041oORZIwN8hyIDArX7akcVki6rglzsVJwZWoDTQKRkO097IhXJWOd0YqtSn0s
Qwcnich3XPZYCNil0/vJx3B6W9dVJEi07Zh66jUQcADg5lYmXJAsd3RHnfTBCBIny5RaOrGTa1RP
EwPSckEUoM2kBHFvIMBdOrvmjRcLAVBcwSY+jTlz3pQih4C5SyDkmaeQ2mfsKlsf7d/k1u8WPO45
Rfr2cN48+eZARHj5AN++9J+vqSCcbsFYpgNQ0wyV/vyPcJb40yCsX3JvJ/wqc5i0W8PzZsCra6Zy
9MGaaWEIVEukq5xL+dKZ2t6Rye6JikRBpfpfYaCOrvZrU30RvJevuDnotMLaL9F7o2Je6KZ8p8YD
3vCIJmwR1083qAaShzy/xmASWeJZcgX5quF+ySTGuEKbdFofRncfWYa2dgX9f/aQmL5WRFkI5dZM
cTPZGaM8ZYS1GX7EcmbjRvg9NBHLiexxxL6XSaBuTP1UK1HEHwskKWjmQvdEpeEjNn6ZToFUeEff
b3QSHfbQUveiciqFwx+d+95/rTFtq74+ZJxavfXiabIySwwxtXNoqDAfMIgBa5CqQzhvnK1Loepa
bpxwIPEl122KJnY+1bzNN6YbceFuOv2OwcsbCL2xtgze6oExBo6tSMotehB89ULh9PD+wh3YpBPP
hdhCcy5+yTRD+1w/s2eLq/+Tbt+w8shhhlb2qcz89j1va50UJffKxa//nTsGqbKOh3kRzgnD4hEx
llVvBR1ZWPYDS63H/4c2dLmF0U12xJupzXAbmsnGGxczC+1U7DwHEARbFSOL3oPrnzbLHVCg3Rpv
Ve8RL5TtXrTeenOUssnE31EjihSbpegczyRs+ERc8VjAu8XWTXcP6ENwN7o/IvPu1rRZtE6Joo0U
TquEJG5oGVza7bg+FXjWVywTPB5srsZMqn2+7Oe+zPpUtNb5jn1vTBHRbPHs3Mu4ndGYnyySkNFm
SR+7vdukOf6cv5W7Y9QOVsYe1B/wWdafbGhS5J++5x1r/ZZqFsYYw/vsJGQzJn2XMS5neQ3Y2ukG
yWWbRBU4SRuUNlgclGesGhok3u1IOrr5b5VtnNLoCDT3gjXCJL1QdnijfshoofOZlr4ilHoBXFSc
/RbMxZoe/JlYjFDYiKVaUy2Rg5WGXj11rstSqEqx5eeMJVB6XKXjZSJALiRcJQRF7qcQno+kgaZn
KnHu7XPQM8NxfV/mhkBOtd+RChiZoLcJ7+Ra8VDkV/B+XWGpt0Zi9LpEx39GuFSqQdN9GjcyielB
YH7asW9Vk4FbskqoTkR3yPveJehN7Zfdi9GrJT0jjo5OCi6FbuB57Z8m5hzU7BJ7WJ7rPC6SacFl
9H372K6iHZQCiH8DYxIbcetdb06ik6iPZPnl4egrT+jDL23q8nydOOZp+Z3FhTPdCt9gTPC1rPGR
zuD9FaXahLUELJSrFmeX+Nq1NotU5cfqJfYUEJMBxTA9K3NaPOq4/8+IFLPOMlMFIu0M4QC70+tY
m7oLy1TMtdbfsssbgjXWady+nz82Jn0yw2mVckyaIlkfA3I9YO10IQVIdzP2cWzyNxdBsFUTLxFD
pSW+hcmNtnNSoiz41i58mmM4A/JpqRIkqwKocVZ11PZxt4GUefvTkK25bV0rAVZ4u9mGOfZMhHap
8O6knt9gtOgH2efWyHyXG8zhpAl5sh2fYKvYaZR/qcGXP8N+g2cbtCChoQijaotsB8EusmNSoz1h
dekcUBDe6WZ/StaxL7d3+4kpSBKaNEKnDKweh1bJWC8FZQcZYFzct2XkB0O/QtOLilyggNe3rbFs
A76k/8bNbny7MaacQb7sz5djNL32lw9ZjyuBWuo9NJlD+GVVhuvZjCRmAuHeA8V9MoGavi05XjCD
R6S8CPj9ujCmqZRpVtNbI3Nfl4OftmG3RtR+f8STevGuWIkuqCV2feMRrFQHcTYxfrgNGaNmE5yv
uZe1/HtvVIstqeZdFTvrZ5PEjDbN4qwOlFKpH7vTL1UYWZk0MWfVJQAlXz7SH/ZD+TQ7Zd5zsPy2
DiS7vfAzJ+72Rp2+eJJKHtQDWgFoRum8mfXViR4Nidx7LXUtIz1tXaa23sot9o2i7nZ43bokfH7A
V1uQo1UEOO+vqZ7nir1n7KdL/p/1zqwt2OYKZPwEXHcQhkQtd7CS4WAAPI3nVDf/w8NyaFmGTlbb
WQHyppfK0PjfJhoRgt5wt6TZHAcmWzFRMXogLzVbx/345BVd4ILISxduvKjQQLjJVSCnNwsr8RyP
ce3LjazHQaU0yHjpDgF/QeJym3/LJaNqpVp/ORtLGV4AQKAc69vAN/3t3UN/Q8uY0EGE82zivRL0
alYx848euqyqXldRs2ZEdapfDSyw4097rEtRLnLVLE19pgxZ1Mo+MP1rpBPZ4f/3tM5MwyKuVnp0
FMXQFXY02zfogdkQYm/GTJ4ZN97azv6bKD0rgkZgFfcheVoJwz4JAX8gR+WPVwvqX+0eTzqpoPji
0uTchaeZ2Dieaus4fUS151ONrYCOJniAHhnSqjWecUEUboCnnWcSN9r+DbEym+c8WccFLmC8OUHb
8n5HaNzfO2pit3fo2b4/N1jkDP+iZRqC88EIvbtl9IicbH8q/G6v7qwc9E1SRKw9KvXAv7fcVeMi
uV7JqfXs/XzNz5czFSt5G5J9oh1MKiAqJsn42uatnEv3rOJDw895T9iFe5bkK3FTkEdSP0kA1aKg
r39MCK6yGQZb/o0IzFP4Y9sXaIBoWEGTk/cyMOW17SJ5CsrXEUnH9/2ku47uTugXCSaHIQHsHINR
zET45jjxbh4wsOUXAa56dIJTeu+/Mb6lvLpou9vosh81gKGOKz8iYN7NE+xwIcpIgVGLqX1Db4YT
KCYMpaKX4nlOWB+P6iAVGjr+8kvxHp+V+Zyt9xYZE4HGknuHtLie8vrXqTSzwI7NblwrXk13te8i
w6pIJh9sfZNalT6gT7xTI3Tf5UugD+p6kcy3EXpV5sG7d3GnjfUqc60qeSlUV752jvhAfZRDZs75
3djoNW3IwKMSx8utcNU+Jir0velM0BctRK4hf/wk/KUdu5LjibCAa+RjiGM5r/958oSk4v0en4Du
KduEtxmrt9O5/9CArufFTpFS2mUOrFm03YB7CuozgzScZpJHQP+bDbQwBnvD3/L0ICn0Xdf5mD+L
XkzLzM22/6UTfT4e+CzEXuwo2NTtb5is1bgp8WkpIR63AIO5zT1soHlRza49UHMexeMeXj0/R6nO
dOfRuzYinUuLdqs8vMROSOPtiCRzFcLzCB5peDPNxL0bo/j+PjxUNTD7eH69E+aT2s35YUI2MWJd
Uj+IkmWtyxrnu5Lush0OaSDOFVvtCl36T3oBgyzdUpqALV8w8lzE1LfpdWZ3JQPMoG0Iu6CHqLeK
j3af00IOXHU0XGPI5ndYnpO9jcuqnWeeyClHZSAZPA7AmIc97zEnUiL8W0URUAm6NWNRQn/z8PGb
Mw6vlQL31S2ZucEm4KUP2oPEXYR04l+a64rZ+F73A2gzON5ikL3use3Sz9diuWGyzuRDgxvkK0AX
8bjZk6qsu6qOfdPEBHaNC/BDagnofDsGxmugeriT/WySjH4nHxCEmirQFIzspw/JYXAcM527NIax
yFO7NFfHQGc1IyQQkOGem+Bwr/DKSvl/pwmjWz89RTP9NgcsbGlF2rI+JtSSvp2OkEDYZZtD/fia
FzLJBkYkYKScQjkLRICjbM26/DzfqxZof7BdL1756rTzXy88LuR75UYGAqKWwQ9MwcveqoRlhw4G
QnCbxvxmc5U8P0jIFLYJYoOZyQGQhyOoUdSXCuZUYuWhy7Zz0RMzYCzxrHv1xHdSAaCYMgzrmZ10
LNTXbga4OoJHpeW91uk0jS0ifLlm226Z1g1KSkdSEY67yzucXcMt2wv26dal2l/isnIptDxXz7Z7
NgjSUdZgYR7cDBi9/kRiMjljNhnGy4nhiwBMoMUFRpumcJxCAXzM0hVw2amTWfYt9hTq14h2uVOu
ESZyvwgYW1aM3Dp9lX8f8fpdjbCMPrr4bZNC+4hIqpOQ71aedGq9HKpKN7R1aNC1UIy4fVtDdGfj
VEzebNbEWaCk9pOeDaYiY3k0WGHD7dy1y7JwWvBS4IyoRhCF1AN/caGxMLl/Wl32OX9gS5/7/T3R
4HUZw4sbKIVXkbOhX6bXHXUlI0hCZlImcWnZhDhTaoKgfgEw5eYpwyoakWDjoUu8ZaE7DLMFvoYK
s9LIIYcx7c/xCxoxDmlu9mHnThQZND6+xgcckPVXQpeqzOpZUrDuRgKWUMrPZTCfLNAnLC08cEOe
D2Hn99W9JVs1sjs/JdbUgeysMkL4nU2dTrzz23nJdoQn4W6RqiHxBJVtOpLrCzEGdl+UNfcTKMXd
h5lUaswHTVcsEfO4anDDK2XNS4SeHexuAhL4fGAI+pMe/JxmZYfg01FpVZvecFmZPtfp4FDXcWNW
Lb7vKpGoYjzA86iEjLGT7NIr9RLGke0zg4sSJq42TlaeS0Sye9HDkltLgBEQS2EsSq8e2dTk9lt/
IFz/ELNhB6UyfsqBqc8oSqks62yVM0RDCSw+mJU9wA4YLZKWGBJyh3Inbci8w4AUgycq2mpsjr3c
Dh/339CvTSAGzOr1ROen7NeRfOP03X9Gqg8TsqVvrxvEGKvFzIHOAIY84iZ8RoLBn91ReDRY2hiC
xaktbAsjqiageP2DP601HpXIWaK23bXcR+rOrYVp27eNv2KYnuPeJkYKV5fHqiKbcE6CVFfgDOOl
VeGrHJgUmREg6hfdknvYnIP66z2LkJuC1mGtID69z1tRFQjjqh1CS2DGWuWEiAoBctlut2u9N4a1
kvl/iJo1Z0QFjS6VUjplj80QE/ngYKSxuDjAwc3Wi5buULPOxCuu+kEvvsgbZqiEm0P9usxBVg9Z
Gt50kiaZEjrBAkkxcw84m+pCo6kLDWoJLofNSKHU8ED32e73T5J44cIdrpSVHimLz1F0Uha7jqm2
XYhsRiwuiNGvfu5RERvfK//Q12Y/MWI9t2bJWyDUsCy19C6UVWZ83V13HKVxWnoW+TuPzvyuO7tP
abUfTMbNlFIdqsWPLyqp4WtWfcZI87oRp81y9M7lI+a3M2XVu9IyMWQMBbrL0el7P6du/gZh3xVU
u7yWNPsdXDduiXMKAS1ZE6FK2SjiLfChhZSx4Zz0SMLpbxV718mPpgAgr2aUwssV8mo/QBUGFF4Z
msqIFHz/hBiBbtC4OreWmdjvaP8Ey/FEqdu+z1WBV24BgGzoRfpaEnLx1dEF5HiiWkCJHvOx2k79
icXrlL1JOaCnVHSQVlxQG+ozUeIkHWBYkzeYVBUfFIjkjGfX52UcEwXa4UC3LDV+gwWuGpoAxPCv
gWwlmVBAtdSjGIwZApmR6oz4EZKN971ixF7WgkUyx7su/HxCMTeN3IyDqNke+1iyB1fYSt0fa61J
yk+3qT2Xm1N8PvUMkOVdOyz59KY8lxfLc9zd5wTEupgqzeYeDbkZoEwCQld3ZmsnQYyGTjIOuGxe
oArBq0M9GT48m+DaNm1UBL5O/D+rAlLt4e63Qtq9J65LABb6DsKluVZ9dSW9EJu3B8AhhmqZ4htk
zOo0a+DDmf839dD7LsMnmw6xF4kGUGfoaqwCGhIA3qbq76MdtdMvZQJ3JHD9jFvwBPGeJsqKjCaF
rlzXJjllwbHD5deNGgp8pOvqY5OBlOUR/3WvhM2hZrvqCxwhQCZ6lz1RyGs8cqtC4dp9eeU5LIqe
IksxwvgJUwDelQS2ArTHQZ7TS/AvCKVYmMVg0+0biiG/XSJFqsAF6WpQb4pZ4/nmZzU6HrZcdoih
JEe969CnakgHNnh9jQKFHc8jzuQNyXx8l0WJTGUQ0yGqKvG+/o1jKWXwTlFBb/Ym7niOnZC5pHBj
h12y7trOz3Mf/Mj1+iO/i1scaHKNopNyMgItQkP/vSgTHu0L+a4q7SVoM/ctK1OGmW6riv0OPGwr
VxSmvdAKy6OH6LdgYlYxd3GAn2bTyCYSAbOVJd6OSwxV3WWEJts5xgltWtDQKVf+Lb3/VlxSUwkD
TwgBsFa740T9zuwiVTVQb8BXlEM0m0a3sD+ndBj+8ZT6I5E7y2JILOGzLq2WBdEqHZytOTCr8MNo
R1xkyl1gOCZqvXWpUVALl1Q5qrimu1OaiOkPeSZ38Kv3B+J86H3uVJKWngs6RqLdWjRj720VkogR
QP2hRo674+4BpTZPEobr4Kr+PcaBTguBP5anmBN6cXJZP6v3a3GbL0J4TsmkgM7vxtH4nW1l519F
1AiIvo6ofP5gaFIcQS1jhCSOEr543RgJSsKPRWWXlhqlrobTOOlT5GLpojQjWbwra0USXiPFot5g
Y1eiHRatpsUZvRbBZ5VrK+yi0mKc1ekIFezXTu+ox5vZsSSLu7pdDLRiAmSGz58iaWkj8ruc8c5c
4m14kZ28emdNg3PwkV9gDGqOXKVjPF01E6qiAOAk2krJEJiA2CGG47J/rtZO4ljG209SbHPsBjkn
Eo8sGMYcpXMr5iq7gE/lUrWPT6iDyxF/19xJLk5Bz6ZZ9y2m6JtGcHvI+01kw6jZQWoficNue5GE
ocd84po+bYkC+zetysoe5U8lwtFA5sNrLTaZU9GrIimlziAMHHL9kKO4u2dy60SR8RfVmK8Okh8u
Y+KLaI+LCnNDu9w+xbK50CJq9q3muemgxbmcxqO9J47Jjmc5+jscm61eVf7zj+sxbkbZ1R66r3lN
G1imBQVyYat+Pq1sPt+j3VieFccbHYCzcFIW/UlUOPcJ9gyI6SQ3jEdW1U6I6muQr7ncorG60QJy
I8fz5bi9Qp1GlJqWV152Iu14Qn2x55WTpMJsXuzu1K02AWlNftmKZsC+Of4r5GwTE1jHUKZeWp6L
vea+5KSm0oH+tnchiodpfTuMW/cgrqjMhqyQhdSm6OhA2crwEwdGP6x5lEf1q3FC1vZ8oQE8m56W
xR4FJnMTCtNoizUjQFhfROf46seEKs/HUH53h1rTC8xYXqxqXHocAV8Xx3Z5Ly8vcTdXHwW6cw/S
Bojp0xI+lOLn5RrXVHrVP+wPYMM0s9q8ne6uHjtIfeFnKC2BAa7RwGDgtqaNtdGP2KSqbq8SKL+I
8IftLhrXm0XrhLs3uWEcvnDhwD6yhJj2jIVa3p4OhRV+4me7hR6pyRSSH4gTmYwgsY76ybe1G8+8
tCrLg3ems7vUpJIxZvS/HXcNVz4AJJCjGrhN/fDCw4fvAhNze634sjp+Q3dJiTo0VohrlBLI/dU1
ccSAYlxwAXtY5iTcfu+QyrQpOf4Gro965rvX9ILZ4Gq/uUGZW+wzQxJS7lp17g+d5wk03HvBj4PB
Q9pDr6npJ4y5jqtGu4ymoT0kpy3jKcWhHQL7utvXrSmbPUDbNhNjQEBm3w5gHyYLdehaTpiZMRNU
HHxX68GkCiEOYaIOXgYKgw0ti12NthowRG2BTv9VdFCyQmDbQ6zC5PTkExzlrfQ8V54LZOdycB+E
VhPC5QhPNxMQzGqZ+U6vm40mmlruooU6HXZFH4ID+midyMkqr6f8Nb7wltqZckhaXbVn/FvLAti1
aBAE26TKdBB1OkuWIdbUv91iM485k3VO8lakQY/5gic706SyKXUWWtHjNppyuR40qTXvMWmJ1qkr
ilS59A6SvIVMmb/iFLmWwHOgyMnDRe6Q9ngmb+4VQOK9GTEuLi1O+EVGTlDvufbLa0/eOqCcdSDk
1HkNnsvHUougNNCevcXek0XPGy8xVbFqCDfvHuwVbp3d5zdZYpn5GuR+VP6qZ1IoZErjHONQ2ndX
EJQ5n+OPj9++vU4inJWCPl2lOsHw7GpS7aeanXaZF9CsKuVk/UAGS6hdO16ipl5Mt/2rVqIbzJs4
5D5XQ7TwoVt7VS+WV+zjxe9uMIVGdvsayrsHT+F0DIzlx9W4lppZnx5jyC7rCjY7Fn4OykYWOT9X
F4nPO+8djp79tH0MlcyD6gfgBVrMtAyGgWCXMNWQgDzrlHFRz7UgXqvoWHHvh+25Ua2wtfMQplH8
vqIPoYw0WB5YBe1Z2OHz0bNQADYFdIyutMrHX2b+ihmUf0FMmujKQiq9xY9oGJqed/ACW3t/xbKs
NE+PJaSPO/GBAYovZl7Sa6m5iV6/eW34OZc5iD3+veQu7zzyzqJs0qlYUWl3Pe72ey4Wi52Y6tqU
rVumt1uSjtLkMP63ClD37767oRRBYxRazO79sV7Vw5pigjWJNY21HzVhwICiQdPx4KzVNlzAEya1
jA0uhxqa4+gqv0uQ9STByT1jVahxrlyQR2K5BO4RPxVOHiY9e6hyl+eCdKv7js3oEgQDD+UUSSbc
UPjF1C5qdpxSeV/azmCbIZKJ3mYlNY3cu7iRE9C4QMiWud8tT4vMvm7HkZc8EpVV7FJIiQL/81gp
BR8mfwaErk+lzm1gALh5Uks75ayqCwMD9X4j1ugCsCB0mjWzdMSEYtMu/yVNQ5MHhHIXsiz6Ys0B
f0Y1IcJ4qpWF5uS6B/yrSOilXrPG5g2QU0KWuFLI/PiYNRVG87u8jjLDTrZq++3LQKZqs5wEf55y
t/6MsDxXwSpAEoHaqy+M9Xo/f2tZeOu/S/wN5Ddk60yzKue9gkZS3hqdGasRENvVEaHl5Pb9kl94
WY1MOq3ipvD5BfpXQA1JLCy5w8YP97or59D2bSCA479+PsS6R8aC6zhmtMzR3O9AeTmXiX+65/nr
L4q/YbwG1aVMrUpo7SFTZwkg0Gdyfji/D6fUH3gJka20ew9Kff9bJGEp1ILhreTjNkJTm5seOL9G
kzwE13RJb+kuUiVuak7m/gicB5SnU3WshtO8P8y4Ji/XBZvn0aZs8DlboRyPahsijZ05ctkwFlKi
FWViG81efJOt1nvdeHOAH76ObpeYAWHpjbcZoAhOB8Me60l1BOngnyy6R6XeuPW6tY2Xuf33h2BJ
5vkxBcWBSMWN75HyjyY3S6q4fCcw6rbl51f+2wjaqr5rGvdLvMfb0FBtUvTH9kvtMq4qPfeiY5kG
iXPw3tSBLH69zMEKR+gpsmxpKLmuaC02z3dBJNkg7mk/QvxYADVmczJ6pfePBX43yjpevlfAT6O5
l4bGxbqAHGyLIqVwXzqO24ZlTmQNUYeMxoeaPL5C+E3TECk8Dt+FVbhryZZS0/kVduVtlIM1GozN
sUkrVzi7kwz7B0PBl0IuCmTp2LUo0wOAWnW4DPUKpSwQvnAW7JiV7tR8VF4kVkfdD4CgiFdEv3ip
urbCy/i7VHmK6djmz2yl701G/+dgiiUx8DS3dS5VR9l79ZjxGX8rjMbC4yOP8Ff0f5kL+22LqdVC
1lgTQ4+LKosq1Rjpm/gm/50nCcm7UcMnY36gHqjYjPdhtc+/hPpHU6P5YmVGQzMja1kTWKOGJcMZ
OjGjCVsJ0rXDlZ/3G12Oykpw8K8bqEP8SVqMaJ/P0YNCPCShceaykjLi9u+RI/68l2p7Yr9/ydre
jtY0o4bYVt3sCz+8xwXMkTEOA1JrDKKF4dI3E3o7WpsF7Ar7XjntWJF7GdK2lpqeevyUroW5mi8/
PUfE1A4k461O6v4n4sv8nGmLk2kJucmFlWWnaVg2nouFdKJL89pmwdKw98w1ENgJxfb30Lz4awZt
YaQqgnfF+Oes+Iyrpiw0Mk8V6KrXdQMvIINBQpnaXfpnGGDb5rJkP4oAgf4ZQLDS0lJjQ/zeLFAs
PwLTRUWCLrspp57yb84O/LnoicdMP96l4bEUsQkWPtCvf79wElC4Oj9+04IHxV4RVIp7cqsA7lP7
uWldXaIV1LYkURDsFd3h39CQtz7hpGTmIUlYGidDs20aEgUO/BHqhHAHHYuW20RHqIc4Z0f+8vj1
vNRzCbfvRwLXCvhzQl/QrUGhiq9DAR8Wfleu4RYKkcPpnqXDlt4W0uJIaDwLSEwJDXjvsVao7zx7
VHwDIjksEUmrI24RNie1tgqml323sUPuLn8o7AcdmyzA406VhkxRejT3eHU3BZ9J3nVkGAwRmZ9W
Zr9B29SRmdrD5+Y8dCmDcT31rt5ZUBw/qCWHBCT+M004irAv5+Zg01AaSX2nuyZ+jgG1MY7l+iBt
bR5rOP0+JhMPPxQEbu4CGRCA/PqSPfkUtQHpSe7+b1avhY9pBAWLISWO56jXRkipMSG+10fvFr9+
hQ+83OfGY1lwTqnQ/9XmG4VYUS8G+Kq+tgzWW1lI7m3NVAGfzO0poaoca0AMansQwJGwsltg+3n5
ZwFgWAJo0xGp9odG6YdIauGaMwm7V9qVV50ZBxBp29v5J081zyi2kmO43xe2PrqUH2M1d2pWzdRQ
tR5vaHQoz5vHh6KrnVr26awf/49Uv9a4XZjQJu/UDHbjEzilQ5rc9df6IY/nrJdISRzaksduUlof
gi6E5ozGWahBVMHCZQzGqu2QPd/7A6ayJGV2xTCKHeoNlb1WDhXpImGXAF6JAcWlgft4zHl+Ly/r
beSEiu+4ShU37Dr1HOXc8EqmZL3DnwZKbisUsyx1gJSIhCnPSqkY4kAXIuMlTUigCnL2PJCaWnSR
Ve2J22d0t4wRFUk0dAwpGfQavK0eEKneiz0SoaQOxUcWij9nWbg9iMI6wDm0ebLng6Tg/PQqYV7m
a+BBM71RvnPlC+CNMM+SgGdH/pA3JVEHsivovcvOLEcEA7UvTZ+JL7+7YONsZ8bRyG3Zdz98Ssux
Sf3gB0ro80eAX5Dhb3UlY+Eq3IbT1vpH0pwsU8KEwWRE2Kc79QMY+2uQ3Mk+OzRYklMvHXO7EpcF
Ab63YxiFPDVeDjTo+JdFyganYWSBSpyQNJTweoioRcT/ZuYhZ9juCY7dlX3K9EsooCQ29sbiF9wu
s/Y5dwc/h3dQIIWloSv062DJ5TFlyWniE3/bsIDg8rB0l1V6yoGFRabaLnetJlg61N+BGeiSqdOW
ReetN80gDkfkXbqg2PNND+jTKOwIwg07iv2JRqXKiMUaWnxccjumPFuX9+4hHqJCUcVPuvnjaiHq
qqiRgvSeqhx/jjfcStzwZeFFOX0lZwOKD6T6hMevxf+dE38W8c7skZdVRysCRyQ/Rlv+p56DIM6E
WoaZSkiOgcz81V45hh/bbT2ddsL+5M28avNvERPMh+LDjnqHgkvhzR5NCMOS4b8Ur8HNFwcd7NRo
l0b5FFg2zNU4rfA2JHE1XSu3RkF4/uOA0gY07lq186q+vhrJtwjBc/cwsDvk/79iOsZR9OYzq8Zm
/Y10rrPTo5pGNCMpdKZmty0jpRiBF7Ey89va89Czetc4N2EH6xQ3JpgWmQBlHo8IiMPA2MTbsrYX
HPXV4Rul4VI7B+ucH3y8/EJxy+XoWgL9v+MR67CpocsRGgxSoxviIdXqk18rOeodS1EE5GcDwTlZ
Ufenj1/zKWXr1gN3o3wfv7neJC+FhiwIh/N7sEzXqccNI2Liqy+jbTAflC5eztFbV4t3jQsLI0S9
2H7SmlMEM7lG7hXshZILchDjFFtm5+BHAu7kcbGJMlDNTL8dveQ+zRdC7UcT+yCD417pHl9UkkiV
GNlZq4B5OQ7kK1U13O12zzwp/y1C3KbPl2Sy+LeOHJudWIyaDY5xYX10DDgjJW/V8qzbk5N2mD0n
J+zcPkCFIuV0u9nab6b7EOJIU/cbsm3929hW0HNYCBGRUspXj0vWpR+BtaH3smKYszMs6OPZqIme
9rCZ39lyJmAwgv7EpsHSGYlSgh82hU3y2xJfFK+93b/tMRa4iwZU35SnAyPIkE+b+8KlD8mKxYe1
aCje/4Rmm152F2vBtgtTaXpC0Ke8cVFdLfIZHS+vZreMx7H1+AOOXupS6jz0xgN1ZEhd64Bn7SDh
QI0fABd20icWumXZSeHJCm90qw6hPwj6bfoeQAswj1Z9vaO/JyS2LIpMUN2jPPK2lsiW0Zwrc3ki
TG7qCIsDeSX5c9RHsM2+VoGkusXRkqJ3BR/mVdw7rEHBDwZLDLCc7OIRDFXTBvfKo/+5Rsyv+m9d
YyZENgZX/Qe/IyKCX/Ps3MI76b2rFUVuzOBuRAcyoE2jpEGzZhHcVkkBwenRwouaHk+Z7FJw8iTI
CmTYxthN3aBOZMg+RGvrKsB5dPg7TRdABRFUJ9s6lCw8ie3IXNhdtVA83CeVD3gyJryK98bCe2NP
MqbY8X71GnjA3Ik9hC7gxniMXJLqMXWqES20MaRfDQVzd5uXl/C/mzIWe3NPPYZYgUI8l8izTvLJ
JY8MCnFtTI5w7ulqkROrqQNoHAcmEeRdox0KR5N/DqWLkCqn5YyUHBAixWiZK3oI1hJZG3A+30j1
PxWmgGePX73gElOvdjXoE0ScbU4bCDnN7FXcFLwUvg2J879OTjXP+cuP+r+Q4B5iWBImvGQ516Vl
L+M7pcvWZ3P61xrXVIOxpuGZIsQoSjwcb0zfI4PlpWL+de963tBsjlcDzuZRuQt5MsDuIjVrbqZp
DtwFIkutBrnJCrobBULJClYJiM3gtjzgRxOgj7Gb1ZYWTFqUosMt2L3htU1PTF88x8Siq8pE7rVN
EBeLqbvoYRTkDX9FfFMtTFOAA1lOdfDjnc04od4np/DqO7Q/8h8xH7vphx0joqQ/sjADHDVtJavm
tWnh0eVenhFCdGyNdEq/DjNSbesGfvGXeYlGGd12IHyGrKPMQrsDVjzBR9hhkq1RKT1Z8NTsmkD1
PZX3/Pj8n19wmutwX4Q7lTH0qXkXZkbR8o9TAmDI8xXtge1bg1TlXfqadvRzTuLympsmjmEFM28x
xHit+xEQO/L3gZcFnDOVM1QgHnGPSB0Hk/1apP4oFOik+bCAEJ5rVlaq40xgyLv4y7VtyyVU3CDj
2RyUpFSFh7MX2sYmIUl1rkfZxll3WduguUWGsUEUj7amJzXkcWhH6hlvfy/8hwdJtQPt8j0ofh4E
Ht6LAXTfUVn+n42a4IboXITJMST7BunsTNpltlTRW9ekyz1TOGfKWznYvIqx84+ryu91lDWEsBnT
fIwpNbORni6iSaoHIReP26lPOmyjBGjBsXc0W8xArh5M7NEppW1QXvLaWuZG3wVzloMaZyLhP6BI
OWRz1ai+WvD4hiFqLn16Rm2ie3VbxPP7LLJYz/mgf8OM3Zsh4j2w9g4YtlfC1HnDdN9+D1LLsIq0
Aq+Dgw7F3ecDm97kSRZlcf/ULQkkoKLWtV3206MrvcNetpYKnym9+TCJ0nQrezJqDgKCYDnvPrfM
U/eUILYZ7jEiEiFhejY3P/9xLtsJMpT5AZtuQP81u9IZ0YPMy03JauJkf9KVr/iUxFSqRUUeEDgh
IiB/eg4y1qyfLKafA9xyfYZw1v9eQ3YxosYn/W/qaKkNG0KI2SYcoa4COhmPyapw41dZnuE760rq
oTMqvpGLcBk4NYMDsaIbBFx0bEnJEJiCPdOqPffCVJul2lyOqJzJACMPrK5/cJQXy9h/tAhavTjF
cQAQgrh13kMueOyKYKW21nWV+cdPkbG5kASY/k84psft6Mu4EI93uy7/f04Cg7SqNYgQ4k329gnZ
1QLEH3vrwaIMb7PnzQ1HWwqVq2ubepd7SZY4puyP20h6GK1KWmpYyO4BLRW+MwLJFUIKZtYpnWXc
bLG5eMKnq/P51lQJugE+nf+uLLgO7VkXDnOb6XRGljmk0RcSF6TQMEKY+nlGpq8zecoVWi0nK5Xo
HCDmjD0gzkMV1DpGuPzMuSkDcsO7IIVLVznM0Po89yiDEbFEJ7OWgwR/sheaJjZVjcdxNAZQ4VAd
k0fD0e43ByZOXwv+RaP/jNyIFpiVlVgtNqLzq/HAfMUW8NtOYLowOrr3iI7i8Hdg7PGSxD4KsOso
yjNRxa76/Mr3PJ0xAj+DY7aUn95ihX5RMRb0hBSwOO1KWuW2Kwx4A2+M30Kz54iAZTy9994ilb3N
DCFZpYJq+yvU7ANJQkgF5BGGiov7aUk3SGqJz8uODE/84Xjkxn3RoX0tKnck8jgYd9jGeFwdcwO8
f/mj26yC52mZAAuA57+6BpI6hdPRxnTuDClrUDhS9P4pUPYE7SjYuzrK1tZ/YU/omxeXju39HQGI
PdrJkFp11/mOgo5DdpfRlg2t/hD59vrfrcRwkBWHKDzlbDfR2IqtuBtpuKixxHXrp0TA9zWTgbAi
H1xlZVO8fbYuQmLKgoQGBqkBmxzmE/6cV3wx+zYw3AyxnLtELMUWnU5kliYPk/8BedyKap2rvR9Z
UOwIlQ6pgxLf+waLSTElHNHEPE6NuDD2AQTLCg2azYZhdhfl/cj5izV+kiDDgtXGm8p5DkRdz6yc
gpvE7q1GicqrYRSOfzaoGRBE+6y7UnaWT50wSo0Rg6n9Q7M4rdl9EyVgPHpqM13VnXSQg3olnW2n
Z5a6cNZqZt5BgvXhGlTjcGR+fJPdl1gQxTTDGbbgvvLgf++eD0S74IIHzSAgciB3MRDjt6OVRnZN
a8ZHR9JinRPlJlMsIf6XwahdNwu3Y4N1D0QkwCpA1lWA4zo+xXGx7dPoWFHm55tiE1fXxgTNL6wr
tf40Ej3C2kri2estz74SFgBAeF767VZvoWbbglNiYOXNhNG4DVoJ/EAvxRqAeO8PCAGMi+unz0RK
sWn9Ok2lRZ00u9gs1aoxGGOqCIFYHffnmTVwrLBoBXBju85WZ4bpoSwFI7aGsYcHX/bnLd/rmMqp
F48K6ov2F0hr2XTeet5/TSMKeFnUQATWCTBVybENJ/5eo931A0zgtylgj7nB278seVPP2OWc6qwJ
BArUx0fmb3dkmg18T3cbZCLmhEhv9N+d2w4wAT0ZhI33zxnoCvjqLepgzOouHWUmPedZKUze4Q38
efVqC8eBBdXqnPPEfFrS0/HWR67eY1Uzd72IZrPjqElhZBgWLHE3TfRrZ5/CrnAO+GqG6rvpgVns
UClQQJiqWzketwilVC3zbKohCetxhmqok4RfsGIZ5PciBJJvpoj+OreY5xylQs8qpCWyvcPvHxZ+
9S1oWMY0Qt5pPrA+3N6F3QPQ/A1Vcd8vdmYYyNrThISF9J3DtrxH72hbOXQaqyxHXlKYmVwuZ3D8
cowtU9xLRmbiyiOP6gShm9gZvvuEqhtti4BAPB/r/0uL5+4v6+P17mxMMYZfCA3DhBgXI+/nJauI
bg4YHExozb+CRpCpZg6GibCgpArq8wBl6CmA1zHAagUjtWmPMCmBKMdM3RT7SR4BswV3s44f5f4z
MYOCX8PVztRxSdes40CQCsfFq5w8eIy5lYDSDFvJ+fFNBpmVLHXhiLUJ1w9Ox8YQSPNUdDJapfgM
FTL/Kza9YROsnzFTOD5Lf5C4new/AeDIzPYiN5QmeeRej0EcpNCWxrat2qus+0cRkeWajBu7so/c
BgVWds/XXU7EHWoQktuoNRfrbzxG6pKFEokW+iYi/RA9LfbE0EanKth6mDtQhxZ93K2AU2K3fsvm
uHBpNoLNKC39TxDcmr1Z2B//xuQ9oyta9y8ae7FDL1q//n+wJKZFIboiqNjOEBaXezQsdWmM01ST
eyTeCzMrKH18IUjLJKov1Sko9xjIr2CJelOc/FV2m1NYWj1pLCbtQPAgxqjkHmaOb+6EI/pxC8lh
ON9Epr5iYfMZoe1V17UNof6bkP3jC8cExz5BKj82Af2jYTIgsFI1UlN1t37jIJKG8ehIhzIfyCFZ
oqIjIODLnTbr70S3qS3MSARPheTMouzC1F1z2jFO/WQDnWmN+O9EGyEMTpMPScmckT0Sn2lp+QNb
2xr+z2uvuq4AxM2+TGSHFHz/23yR7C+zn68aXJiTRUx+66PrWVL7iytDTWC8YtbKYoCpFBIqEhqO
EU196wjGqyGgiH4B2QlkhKb+CJEdBwC+nnXI7uLEM+ZT7LtXq9h10YbAcByg7sNHz/81erqRWFex
HfXvNnufV5VZBRVTJNUh3eKou9rhtH34rsWpjmBTgMcQQ9Y/U15Ql+CPMQOgEosOWTYy5k+vLPL3
eqnI9U5ISXYkP8RGzj6jmxs9rYUyaz4M9e0RvKiXYHJ19pTbNIq/DJK/IDIy4nC+RmKwOv3D8hyo
jqDc3Gw6ChQVbuTZijC9AeIqAizfOABfSJxPouWn6YUAVVUUFuvwa+wdkjTi/wQqDAnIQqajK6Hl
sfiwVE49EFqUOw0t+1LXX/dBmDGMUyUqEZmvyRGtzERFbD7qfNY6cN4mW86ypvkbnOqCUFd6HSmx
QQf2nOsu5lStsA5z5PQtISQiXATdxU4iL9KuIzSiSM+eV95xyy8Uof6zpwkwUYc+yweKB4v6Qlzn
+8Qdqzd/VJMZYy7S6SfLHhJ0e6EWnLEjMogtVNwLb5QF1c0or+XKmlGISk9e1R2WPsOuMmIFCPQM
tHRMAPgTlyGXbQ2EJ3YPgsgKYKkA8OncjGn6EWv5pylBz3p+b4GFuqQb2aifqOVmfZ+HJgDtIub5
AkoJy6kr0q5MAs8k2pYqG9Kk0/T3oiU6pZonUEQ9lefsvuYK9+vU4ZrQbFc5IKejXlpYcjWk42Ws
B1gLmi4hPqAa9NoXsCf5DYPQ8f34JsXif/AuybP4PiAgHBhTTW5x7AvdiivuX8IvJHPqhpiMkY1D
clZU/2AH4lbsntpCDlRx0byxy4FwupfZTGiM8VE0OxMEUPh3MY6JVwfmVr7ePe8cUkSNh0R8f7RZ
1EdKfSI9F2BW/TnH8vwQonSWaUNoMk3YLQtVtntXhhoi2HZAEaog4c0aPnibmS+nEVZmxUx1CmHC
2M/G3RpVG26zGtchUH+Ytk5lLX8hECD6/TkkcL+Qot+8QoabmP4Kz4mLeUIDv21f5iZb46ZQdsvo
DUKhs0bxBAq6n+JwulkDxpwrQXFQ/IdKmorcQECcAHdI3YNs0q1CKiQL0Uo+qpLsaV5EhVICVH3d
DON47sxsHEXT+Ll2mARah6+snXVVv+sP30HDa4jLEin5OLyh4ESZj3R0Zgp/CK8MXPi3aq3w9los
u31OycV3/3U1jdWSkqHnrkHRg3Tmqkh5c4utRL4SFkyxbg1dVHZSWxvZllrdUjtOG7BW/2urUt4X
CzyCj9Q5yDH9tRkdB5Tv36odJU5Zlkxhy7Z7bd1/mG4IlrCjRR7SmSggG8FLu06sZU+wl/7mA6l4
FftBaSMfQYPSNsi6LahGF1dSEmC9Dr87qLXEZQkxeaNhFnio5LNkOlVw7laBskctpuyYbzGUPAA3
2WIh5pAat40HZCNjeRCzakNTvdxR3QZCqA/+rMzy0lxmnti95npN5Rua9cAoHdXsysOkqKafRf6Z
2X89vX5GMuQF5irKg7ZJrI6Br7mPl5QJnpVSvOi9FAYjlh5x4ns3rFuHnfZdrHGYwAaUc3sEPAKT
N7Dn1T3sc5o722d5c6IJ+ai36zOhdX66LMoGPuj04dFUrVJ1KwTbcahhSMCQlg+1elTyZr2Hg+1n
gC9OSLiOgqjhQCwveJXSUqDefkMIRVrgiTcWNUa7ShMdHNfGAOzxyojjUgqbapluD/6XqHY/x7RC
g6laWOeb4B9lw5PRVEo6/Rn0hXU0eIhljdr4+b3oe01fNTqa1R1+8ulqiCROkQoRA8AHWQwyC5mR
qxPDQUw0sNP+92PueFrvLsMnM+Lxrp3isLGow93Gl+GsGAwCoWog+anh44L043hpdWwnlkpIk0rs
i1BeHoYE6FPaz2iiO0LyQfbjL/AFSMfMaS7P3Z5ZsLV8V4ICZXjuSCi2sNwMNTz7iCCIK7yP4sqd
suXpLcV45ArD1Dfm0oDc2VkhELNBvlMz+uMNrbPd0rrGFFPbBOVSRvUet17xh5Hh8Vr1KXpng6mK
miVVc/hgDW+OP8eItD2ixMtHL9Sqv/JojdNfPzEVbj2oYT3ABpeQZ7C/NsvVmRh/Q6DWVr2inmaj
rSX4HMijs81yevaRT0KPmA+IZYF7R/Om3YzKab/08yvPGbB3yQRqokGCxibBHE8PFYWjB+cAjwda
782bwpjzqUzmixiqHBQdngs4RCLiTaaiBs4D6eEW9lpfl0fvqydtOimjztLjrH/g1dE/ENFvPZ8N
PauudKIOLgGajMqPv0Rrn4wFv3W+CCN4znofIxjN7fzcRMXzB0Azv2//PEl2qyfnxxhKKYLY519j
9HxdiPs/UH0LJ4+9JxpgMw/pNydqoqhvcPI1v+pt58eX5k2wRrhHDa03JNwYlXgJ0ODEXj5oUC/w
wlv5VqobQ5Rf0bronBapF9MNwHKeMiDdynf7x45EOYKEiT11iJkNez/ue8/2EZZ+ZPuiPbFRax74
5f5EV1GbFsmc2+PDC1wk2RaphWlWmo2Ur97iSqBsSfevWhaNcG7C8wVG4ogNJ+fNCoiTjS64LRqO
iVx8S64f8DgSZ3a9AImZLChiwRcOSSV6D6LJHz5CyDjPaVRP7YFIEtGr+kt91WDoMAgP6+7W8GCt
JlxR5ThJLHOGuan/+6SIjvdT6ne72VxnU2A2Bgr4WK7ve7fbIkCOTP0f2JIloRM7MdCiK5JCnsRC
+h3mrpMVTl3/Zy3Me5VQvHk+mN0S/+eurehMJRikKsP6XITxm9Sq/AOUii2REjfm/16cGv3WbSIo
oTUkh3GFSDCf+0H6rZvTCt1ETMC3NzC38gmi/AO/mSE/We5qLQ4afPBUKzPiKIcrK3MNQcUFCDBm
PBkysz0EilcHIxdxJ4cuDrXgnmH88bm8ORIRrgBo52WDPsqM7GVYG6yFpdCtSj+EUaLHDngQcjMv
HMyUOt0a4kckJXf+5PYJ3/qK0Xrcal+yVeqFAh0BSRbnn3hocj0+YuPymuA3USXk8Jlfr94J0Qdh
S6k5gW2hQfknKZuqnI6UTIRKzYmXvv/mU3S5lKgbibDJfDbMzgAxaiKqdoNIPGQ1JuJ9pkwLOdIo
lK4MCraxOiks5+6gYRMrsOUuZefl4w/ctcuT+Z4KBZUZbZWzIOM74RI2S/+rsYKn0ET2Zhbu12k6
6gDCLopElZWlLYBekerteHQszb3QAo3h0HTbAirkopVnkkjmNyemehPMHOLDZvHvs/QeHowBokgp
yJyfc/VIz8ElaTh9macgpmo4sk2dtEf36Z2uV02K4IAb1i9V2h8lypYeMTboHhsrvpxvfH3YDaIK
PiFki0HsjD/WmPpoLHpkNFOYA2UYIpX1GZOtKCVIvlWpFtXlOcNNXkkSzl88o0U48Db4zqJbjd/j
pD4+ptHtYuz7/YSpPIrA1kiPrGdtSYf3i93poGBWUZ2+nEqwpMVaT1eaw3TjgGX/VeirPKNiEoQt
CxdUEwdrOcmTBpCdF+rQbTQCu3eThfkrT9hk/Gkdo3tUokYzQwr6OKIyPGBpA35mfBbhChWUQQwW
c+X93gTk5UDTL83Qrnfd+dBHWnOean9knVmf3VN1fyDS+13BMVleqoGt0K4ffpzcl8FL+bRv59PP
fEckrXCGGPY8k/w8KQJ/Mh5GA1asmLxqVGY8urC8EqnZ/H6iK2QfZiYOYIUTgsk5ruJlK3++qqbI
47CfaSjHQw/7obLugzMHWy3HNr/NlIghEPFDrnFbb1Ob4a3iouKGGV2Q1W84iboY77Q6Roxe401i
qvtVzBFr/gjTB9JKtnLIL/McphJFG+MXgyOduqr6zJA/bfYFnh0oJjkLa68S1aQ6tMjrP4hH0lAR
J1V2M3lhj+DKsxdnP7lDf8bX35llJCrqQewqLjoM9N+U9I9o5NOUqAwWUEHHqXArlOuJ6tOIZTrl
6EqTdlc98uh1Iiicl1FgRTZ/QdKmBw1f/W54uZ7vMFcspkku8lly6b3CgFcpE8NY1gt4WNYMPtSU
kboEf1xkDPzr8k9fVmI81PDSIAuf91I3uzuEPAeDWVkrZnUig/P6XZBIoJVn3L6mntnejPgQeSYc
i1ljVqn3ldmi1/3jSrrfLa7elBcXbXkz5vlAa9g+xLiV7OQObzHqwE2z7JBDkNfMAJ2DVLUFyeW/
z0lWFufK6VtcZ9YVrO6HkME6GlEwGvKiFlmIylZcsy4j3F8meF2v9St3Oz1KsQUMHBcP3IRHOeca
j+n0k8CvHYAJ90wTXuAXVJoJT8mW+Z9YlTdRyTp0Jml2kekuAHarkkmFIP0D+dJT1BdFrFS8c16v
5XnJajrzsG9udH1FFNKfAJJbXR9uxHtCaQcEkn+fXd7/WlNplGEy0YPV+y2jOPS2m8hzvpecVXfm
4UE5Nm92pSv5Bdm3onNKEuv0ATmYz7wQM9HAOI7eSLA80snlLMGZOBjqrHTE9jI30N6mOweSsd5u
4cihL65NEYUo3PgYteAY34CGTvLUoqhxDRSsqggaw0KeVkwitICpAl/XlulC7uYSF5bUqZtQqt3c
6r52WNZdMJbll6lXX49ShyO77I/SZHBmCKfmqgYU74v6cpndzQfYflpY6ZerV1/hYglcQXA1SkoG
4TcbPHvReBWjiUHDo4Eqet7VJkeA8+aTRnzz6dQtSSol7V+CvW3u/kPmezmrVQDJssm9N/z6lKYs
11mrXTu/VZLsPOQO8BEM4MOv2+1Rve0Vt8EjUn2iwk24fnuMbtasJBVRrNqcCIGn41PRjUyH/6lY
donbHBxeJN5EfbdTfzY1CD7GDccPBkUyE7VmHiceJfDuQOWRjTJE5YViwJ4glgQYIjjDKJxFXPSQ
91gRGUG9vlUevFOFihSpfwhPoyh0qF5vngyAWwF0F3IblTvC7VtP2AgfVDf+sLwzOcGjRPCDXQ56
eK4+9U/rze/XVgcdMlXx+sovd++NqbnCDWOwRM4waoy06wIdZ1/2MxvMZ5knf7aryLBMV6mpaT9G
rGsDVTITdfAg/Zlg7G9SBrFUv1HGxI3qj2uNEEWaP8BObTJ8BCc0TAZFFEpNpxou0EqA7ERapLLc
H3M3SYc54DvcXFo9d0xMwN8f6eBCWGTRoS/Sb17vCsqnIe37k5cLWbcpo3ydTfJcrl1dlP0X1Yer
Z9iLwHwAiuEgInkmkqb7yxXRwUSIYBEFvtfGZ4+71ktvFGmW4JnCvaETx1+947cTFgOGAK1p915j
JQWK4FXTTKFsFJ3Mu3UnKxMXzTYjtgyPN57b9pKdFEurwgzhCuiRaqv5SNNoUnkFuSv8D7bjS8jV
yUzNvYem64Ln6GpjfSRaS/M/sKnSNMrx0NV6L4b7SJ/pAqaeyO4VeqowxoIXkuc15zjcbYVBKW38
O+5nSakIUK7BcjncnpEWH+3Vvobd/fmaxfqWX7scPkA93wkLaRVTmoGjenF57mHzL4nMcKE7dz+X
KCXfCmiUaVH/s2v2oyV0lc4gjybEDOJZy/ecblT+4v3qNvbdp9lGA02xkw2GWT0lN/OK106lDAS0
fywDJ+l/heeqw8cXeFDBvwPkMptBbbc8/nwotm7gdfA3qs5l1ILvEQms83M+57yOC32avEOmuHea
2MfHCOAqfFOO4EKRQ3aeErSmkOI6WrpunItLgFfI27rE1eYunsJ65GhKSmcKNjwemn+C7wiN3fNN
S3nGMRDZV9NMhek/RygsvFYleuXrcwSIfgmXEw7E+zdah7iOMTKcJ0xHTSw16eO9kRNoV8qCrLmt
6NeQgYjiRcVrQbSAvwnZTSIrD5E9qLxx1gHo7SDl4kUhhH3NKKE4V43cKAn8xIQdWoh9GWPH9awA
0RoKe9Os1SGO/7NQ04/aeb5JGqmr73ORkhApm6aw7GMcA7+PTykTviIp4f657s/44MBz45N1K3Ku
bgtKbiF5Iot3LDbdceGrCPAuRszo70RlJjUm/LmXdcwLj2BWQxlKMKUH/EzIq6wSbp0ypwznfdSM
9p2DA2H22IPS5FaT0l/SVuK1LPY9QHAm8xDbfXvtlnEGSROapI7G/7ugwK6nryX83N8PNpZDcQL8
GskrynIJkZ0ZlYrLCry4KPs3Vnw8tOoQ1rlrsR6Rz9QO0zZZykm6rTyDzVYsdDcb/QrC3fSu34vg
+qDsV3cq0D23NPv8pDDKNmo1LQdYwhw/v9yzOnXW7C8UISlRBRaXrAXh/EF6IZ06tB4TWPnCR8cQ
VSuqu8jAEBvo8d/I+Cq59HN/DpUrZ1unYoOD+V4gfoCLerzxEtbSVc67m1jlBspSVuoxzBPRWDne
dp2YCLFm0rEsv1e9yD4batJUb2iQjxfice2hmViRKuV9PEnGs0QM8RVvDEQRR5sKCVv9E2eV+0Q3
Yq2RSh3DBql4uRsAg7a/6wCzmJWKwwn9Golt2XS8Y+rLHJS6eysjpDPWWDoA652gRw/aSsbulWGu
dlPfsKussAa88y+BaE0rgoPLfg8prqRUAMF1kB5BKBkvtQpqniqZ+f1yok/QzGYQ0CZAtfejFSOH
WdVAOjLViO+tufvm/k3mNi4vZGDqffT5O46apzw7kIrNEHSlNPci1kk5nrlmLPAJLSvhKvUJKfUJ
ot6PpNbkR23syodU/m/BRQBdRc2Yqpar/pYcF1hsbF25ke/bdLhsnNv7ota8Q+LlPQcYjqsLVRnp
RAfMs1i5scA8nk2BLYfPJiI2juBlIR8a5+rl+iMT9XGdW6w4iMMYZMDnDCXRv/eWGThjchn5ANDT
aZLxU9oWnIj5hC21CNv2/bkpWit5uwQv9bXXl60aG+2yztPxmV2LA15iiy81ItQ5i2OvMmi0mG0z
DSNvNFMquw0i9BLPyN3jYr+EFoQ+juYDsG0D8CDMYdpYZ474lj8dH8XYHVMkI9tglVz+oW5tSGHs
NL9GhV8e1CWXmLWs0ke1JmPmDqqIY8aVoQMoO6fLtHpiLnCyyvnarEDQaHvnHm4121biyacRY9xh
J1XKFJ6QDMhAgVJ6LiVXZob5riQMZcvkbLy2s3D3GyMZ7x33Sgny/wK+OSGzHX7X9BXrK5HT9CZQ
0XAZPfpQs0Al4RRjKuCmzwUkfGWHQBSJDR3oYvuwpiKJqCR4tuKYVhhzTthAqozV33j2McjMRPQW
dQPAiAlFQjWSbFFEUoSGiBaRBzGbTD2PItfKSb3eifT5lCZk2OJdXSCtgSqS3iOKLBh804vFuCmB
KTGie92dHU74SCdiUtbBCYTpIEckUpxAxnRh/7iWwTBE/qK7x1gzEFKvCebXFeUY+PfkaattbUZ/
U2b0qwsc68YOgC1l348xa7SGKJArraqKOZdzRnjnWYbL5C7Y3oCoLtC4HfIr9NY/qZrElDpEBNUI
RrOwMHrMTXCIQbUf2rDMmS6q9e4wyDjtc4Bp58ektwOkaLwpa2pmeNgb//fNC2Pw6F31tNKiQGXb
6wOEtMwQBNaY0ZMYtMu0z4U1jNeP+sFYW9pgCkJkVtYqMkBXj8IS1+7ryYwBez5lofbyZuGq6gH8
f4vxwBpsLYlX+B3dtBZrw+ZTYlXD5TZG0fHAmn+ufkV0OqUa1O582U9tw8IyXBEesmxEFc11D/pF
CfUxn9bd8r7CVGZXTXb5o9ubtDAmjD6vZESDZvAAAnreaXi/MTkp0LBuj2foEU2JxN/0K7FhTEfL
bCMPTDrFuj/IvFNCYoSUF+HEH9S8wcUTzz0PuJ7Kr8Tc8KWYC6E700DjzMqa/vTu0uilUaWZ/QAE
4FUym/Qz6Fm/vIpkN+mOVtr42sO01t8A+52lu6KTviTgzf304DuwNkrcijdDielRTasJyQm636r6
E/7v8YF+uoYsGE5k84sc2chTqYvS+dgBCRckhffB3GRv0V4xxB7hxmGin67cH7opdJPSgJMNR86m
08UU22pby+leqbQG0O0Jla+tsmB5TZvEmASBjOKbpumvv6s6KVJ7vXmFKbJmXgBtUwm/Z2dWC5lS
qHmQ6pLU7lC+ilPn2itRUaMFjmfcX+J/9OBANjXw9EXpbwkBvfo51X6/RmO/nTGYb+HVZz53OC9i
xypP5vVO9p8q0b5Z1A3vvBErQf6yEanTAYjT6hW+FQbZGp4as1n+BKznfwk+IfDNr9qNDIzIsGD3
UDJ7Sj7UqmQtId4+VKo2g5RAWlzI+zWNOKkPMpNAMQxccrCJy2+k7cidNClmxpKyWL5UO6k95Lur
a/sed1oU7M+j4Vp4V73GJ3O/1PkAKf7dwwywa/MQPeiitIaVrbu4HiU6Cxm/OBEWkezPDmo8gmHW
CLWV22M2ahIdbbqe34h/4cp4NvKNSl/t99ijgMbIqj6qBuEtzb66CIdJ5Sy4bRw+8mFiBdfPT2Jd
dxbid8Iv0Fg2u3d+7OxbISOvY33Aj4Zzsu9DsIlzQeh9FQ5IB6XwEa3A4kJ4aBZVXD36UIo3DkE/
uWSvkc2kN76A4kGWR7iH5Cq8mdJlK/OWutfhsNpz0HYQ7bQbGBB5L0vACvj7JjHdq9xZ2/qq1qew
R4ZiyUcIpMBIDbgpekQo+fOZp00zfjApOkMIg3qQrXcMi19qod2cVnri4NCU/ULw8T8lbj5K/Acu
2BRFu6jD3aqmlA5C0lAXUmREqveKl6sOZ7tb9TXzAzCq8A7D40WT/OpRqEzlI9T2Y1rhICBmJPY0
zwGULpdnLkJht/DDXQByDHIJRviuh/Kz9TYRgImzVnMhDZ/al+wljd/ai8hO0E0pGIONm4fxsWYi
LnfKAF5z0vaZ6TnQRgfW8tlCAlajAGgiw8OlRStKXQE4qzXmzuiWcEJFtA2zfkF5KVwlY57QwgO8
yni72eHQv6+8/1eeTb3dSUGmzrmtkZEOstLJuFPrNhacTU3lvkFlY2pr2C1tIzcCx0T49ixDTC8G
jLt4cYa3o9z1n5mkZznhgzaPaSmYZn077cBt/Pz6FZFY1VTnh0Ekr+Z/rztknH66O6DAdlI6RkiA
Qgp+T/cuSKoh5j0/lKw4CpRTRHsqcrD5i+aO24VDCu8NJYn4SQEJyU4IuniroZhyUU/b3rUXTMkN
RhJNpvt/Bpc+49UY9JDIDRYdSnP1xXX5SWvEN3RWxWHjz9ATIp8Lf0QJvwz/iBQc3g5S2+YLNjH1
ZU5bM4Cjl1Nwl+fb5V8Y7DQPezu/jVaaIGn+FQIomqrx8EwMVyk6t7n6zGsgxoxci11lUluBn6wE
AQKOTv7cj2l0zYy0qtZQG1yb5h78MnFNd4zEjvD7kBxDU3d0CAB0qQK2DNAQ+Eq5pV1AslTvNraP
JwOV5MiGLSyDRKknH71Gr1cs0CW7hH8aYDiUu14VD4kYla9hJmCctal1Dj8BAU1c0LS0eai/ww8w
mSwqa0/FkBozDSU3BUBUUxofLFaVKB/oruaSs54j2v1xc+sEm8EF4WQDIwxdycWnvuNLjVyocsTB
hwHTO4nkjEsBj7nLhHCXNSjzimWIXkGS39ECguXcYIcW4iN6lGRjvqga4KW+BlylkaNWZ/1cGTWw
GPBfL7dt/ov7VgzXzEyZo4D4LM0L+3k1wmNq74V9s5tu34BsuCSjev7LiLFHII4sDlSrYQnSIgV/
hzOCxBFIQ51QcCtuMTnsmRIvgC3FvJL4pDa2Q3M35Lh7lNge7mxo5bJp1v3N7UsXnHcwO6LzR0bg
pTAN2/MMv/J+Ax9BRPeW0aP1KLh8XRZKWKmihgtqmOWrAc8OICGD5sbi1AHp2qX7pZWf8TtP9gNE
qbW9sCm2vLek0JGh7wnqWgxoO5yzujbnMHHJ5laVSZ2s/U0L6ISY5PNtgm2khQLTsiOpdX6RkAUJ
WNbSd+HoRAhjHjz2rEbkVeWXQg/7kSp8+VUqDY6nqnXeOycZ+/gk7sum0tyl40FInHFsTOa/M2xr
IqBjvqI82k404IvQQmMGnteOaqNrkODXv8eD5qZTnsfiU1cfIm4B0Bxa9r4ggYzVdqsrWzFLa7C2
X1vQ+r6VH7zIW/mRU8+oNgmL2mYU94W9oo/25gucex3ZmAv6UqJc58a91/vmD4qOwW91GwtrpKkh
o/y4k3NUaHwx1PZnLg0jWgNUwOj4qyVrtyLVaCj48p5VUr4iMZffo6tP8Q1fcIhxeO3pl/Co4qny
k7O79a48ZBHnloEWfD1PWHoYBD/vFl3ElbDDflpbN5SgyyPpWK1s2dezf8mkVbvQPPaytNMMUVgN
tU2Csl80wJMJcBK5DibA+JCwdA6SxeF3Rrk2V55xZu9z5Z0/d/gs3Te4iRHXQlITiZI4OOLgdaxI
/apKq9vCZ2OEt+aKG/lNIpnFwiVTOTlv3bOsp5M5k+1uvsfi+P2oq9E4ACcT6w2ur2g7XdSXkllk
7A+bU5X+Kgua7sOr7Kon35AgH+ZfvvI8k1KWYc6CVouvaQE3QKrVTsgrTE766V/1zFpt4TIvSpjG
ImKOuE+bu+/wQtJuZQ/fNldRPO9VyYQBaR7NUDS89bxXl8WHYhbOrVcSlfOma6wPHcS392iErRvG
17monNA4ru0HI3wjXNV3NojFBgUL6RtxeZabl9qWH3fLXfH7HPWyOwX8wYVwEKh1kKBcevGu7Iiw
/o3gozdZ0fCaVWjonxKQOzR3eu4e4Fin/OAwmjEZZJq5Q0G9rPEm1bx1JjAtDiBRjSOKkpCyBr5y
gm9CkbiVwR9scpFpEQwUDYRWA9H83XB8M7YZncfZAFv8DFu0uteeFCa35QOybHgWF2oeMSKDSY36
n52PkWxP80jrS8Nm/58NIX6qx3MN8V8ydcaitG6TrCZjJhXfrPFnTBGQzinbm/nQrtGvRLXdgG/e
K9Pj8Mb/dQfYGjOe+WJ5rwR4IfyDB/nrccBeqCYaih4tzR6THC9R0EAAkhFVqwiLD8/4/VOpU9iO
LlZJfdpK/4cHktmPR7Sdn+mgrrSEzPC+EYv/2UO36QglpvtjgZWLrZ517uaGUFMqVzgPkg9IQA8A
zkisNYh7+YHBMPEEZGmhaWbvT4L3ECx4sAUqEFFr0oWUVHlk2kSeVRC2HN+x/9TWBZ7xzRYW67EG
Vnw2LMzJjUereTpUKIwlx4I0SS9qtAy6eVJowpyLjme4zWOvbY8JCn6nfgnBaZI9roRAy6mEBIjS
A4Jrn4iiRQ1dY54HYk5brCuw7OWAuEIb9cMlqEWIaFR0j0oUln4PGp9e6xvISUGgNsIQZWo4he39
AyS2GZuA4aBYNHdryEolvjJmgRgNYWQlycH0HDSAW7o6ZZUT1uon4X3SlFl06S1vRqc7FsBYAnf8
Y8h8rB4xYMZHmmoOxB6we96J0YK+iGCnMC8pDcAgVNMSHoCXd1NS3JIwnNi7s4Rov6ve6hHp+/37
0+FSFDvf9xP0ll38ZSRD0Wz0l3HlrAz9SMtog9UTPJNcTdH88eevY3bOICTxEm78y8AR5PL3O6E3
KD4fdE07u1nfCaJlX4/dedQ8NP53WZvWbOp73Xd+I/b4s5JElxX+A0dOoU1Bf0VHV57S62UMSazH
OLfiYI8u5+jGDQ/iAlb/Uu2WfQvGXlr00FKU+SriCUgRdkGaXQIKDvrdcloH+eoAb/i+5YsCTjOL
tRWa32IlCKaERHs0sgrxK2rfCorJCuITTUAZvDT8PziQ+KY4t+ZN4HDHQPLsGDgi4TUEMAJhytu9
LLCEJLtY/PUfVb4Ki3/rqjN+C89nNMm3gqoWC9PjUaWHGwxH6GlRPqP4rAPkfeye8HmoA1y57qop
hfwlo2A46F1XUttlC15tW141wYrUPl3vXN9Yu31/BPsqb7ZV/ktB7aZBDio7CahxVUilr5JKkgCG
AiokGGyhXp1w2Uuo/Qd2J0+j9gWOoox986z/vPkQGRrhCp2xUZrkxP5mKtMKX8txp9+T64mHc/J2
z3i71OOCJw4hkrFKk5i1KWPj+bWxVWuLm0BsY2Iy1zghMpxRsrfg19udslAEUGRT/dtW4FODjM7k
e/H0UNVAcgrzb4OWQs51jp9P7f0vAhPR57g78zOrr5/vuj0YfHN+GwQeD8FtFZCs1PG9+bo8f7Ik
N+dRXFBNaj5piYkbWF/KoT/cLnmMif+eB5u7vm2eQ/6wmEekZulT8M13PVbt0h4HJ/I2TiqlwbvJ
WGKtvHSFGIaPF9Gq8yFZrWMIfUwnCTECux3QSROIeGMVrcH0Acwz4pklfNq2lulMmGYtlG9Uiky8
yKq4HuDGZVUDJmw3YteYhQt5bMOyMsv2AhL7sUE/aqwYnce28pqzy/TUDdQk6wcGFgpWOJaxJxTu
6HDgtd1WrQo0GdoJD3Qmj6axx9xHmegG1KvRgypNRIzX+Gb9l28npOtbxNKaII83kl03yUrQranj
NhdqhjM+lshOr/fO2XLJ2PksCLcoM1g548ZVgGIVL0vHwLI4eySaVZBGHthy1zsi1i0yazYQRZKU
u9KpxkJFKlAPwbUCLA9vwMlDp/SUu3BAommJhr3oDD3+N1vlNXnmz9e3ccpvvO9YuU6DqJL/wMFB
R3T6MmHBKm94pXosm3eEVP8+DVHoQV6Pvec5dzjP56BOsXAheugdbw0WzC9ePmYte45bLyJC+Uz8
At2d9XiTKV01AkqwVT16SGoxzreAkUO6sEJkulkYz2M0f9W6tK8NbRjpjjXLjcBkk/mPE2EK8v4s
m9dmSuZVetf+D4EYTMl9Hr+zDQQH2/JgW8PZuyE9mSIp9ppef6BJJcGKT+p+/JWMRUA4rztgFdzL
jo6rTjfdba2vuOFfnDMezEhxtFqBrHog0evn2brthg8LdYNwZjJScbT/Lo+EVMxjbm+GyWMu4ioV
LAKVXSA4Qtol3dPkgwqVFArXHUDMtMZpPzx4dUPEG2oUpDniBn+eUtBdAG2GdWJo5sf8OwlneZEY
vm+6I9ri+Fyrq6mWw9ZcuI6B/yPlOb0gKp4lmVNZshvijyj3Pp6RgM5320O2kQBVoMoaDBYCEDRI
MiYQUP06weYgItfDljaArkXMFJO2s/gdjrgpzGVhc2UMd/shpzwsDcrL7X6pL/BcC5uOmEuNoZA0
CNxOdifOw1RZHVXcNEPynrk/osnCdwBdgJiFU2HtYlSA7UncdHdcyZ6VorJ9xqddkTnrg0SQKCfM
mW5LKggnjshDbVIQifuxteWl4SlPdjefFlOG8n9OyHzgQ8vxXP5OWzarEtOs1L+0iDnHtqsnn2BG
ohL+sjUCXokD34cg8/BtU4QACYzXeY5eiFDL5Z/LIxOG9lXbQn+u9zQDk1iBg4Cv/a9j8K4HA2jM
P2TsuRjJ9fruHgPhD0ymHU+Cq8FBqc8lO8Aww4YJScUH9l0FDz9JqAu+COskCgd4nCKNFPd4KvIi
TX/DEb0KaRg4JBPr2WLrquT4pZVBlRrirlyJOcoaFUxfebHO3ZurrljxVKWlDVC1Mu+Q5ArvG353
cO89GiVhmprbWMUUwHCsEZgDJzBy8OqMJcnsjHgWYWPXgdNmoydZdaqwtCKIN8yCKiEkhJQKGMC4
beKRaapcizpRX+f06Gq27h5HCaSy/mm6onPUiDSZSZfEqHXqjRI8NETezr8QrZuL16CXjY2KASbV
iklk6BWUqycyNbWEaLVSgPbfutZEoOamWl2hdxT8S+tlHhBxVRJg3od4yevzBHbF5UGX7P8Qndpk
Zz4qcvL6DEWSZp+Fyt8sDhwc6vuni5F2TPSVXmZPk+a3il0EOogpWD8dzPIDmymF8URqu5RTVbru
nf21/9I6TQJwmwytCBwjNhzomCZEOfMY2vkkM0DdpeP28zRBW0us2ZbWRmLv9dAzgNpdLMJu+Mlb
FUXazGiXTwJkyRFEFEqEZvszD0lBeEb3509OO3ZTifQKTyHgr1Hrg2aAXTngZjPnEsYzQbNHkQDa
nlZrDGQfVOYg/qcynCrZ/EgC7f9GTj/ibj7uQ+AJuPZ166xX0LxsFdm/OxnReLBacQbcZXrReaqA
giaM1L6HOTBtTTF/XsZgW7Ie6otU6YHD6UPWquNAs+avc83usEfowjHig7hPR0cH3FdBCIbwSgmv
9yThoxCIiMMyr4jeciv9BtdMyaXCkVYBg1vOH9aJoC14MklPdCxrYrDDzNHEzsjWymLYmvXOChlY
JiKBFqB9JTPtsPnMjYI+9WRSN0PKcrf0NAnaoxriz3vf+yJOp2K5+L9mB8fw2mA8DMYsAtAaiK/9
qKQoNxYAahYP8qUKKF/HG9vP0kCbhAFT2Kak26ykT6a040kzZmmvm1G2WVFlVmtzaJqwUz9dacse
4TKrm1EUtjChPrYbriko74529Y69gfM/kiyMJKQBFT10aCCjusNgnRyjYqtPZlFx+qAGmi+daJsf
OJBiuKDwOreXZvRfwIseqchGMNcfqQdPW/RNB4XkBMyD6wIdknWX4twi6NimUlRjM3kSlMnv+iuN
CdAnsndRIe75BSO6h+vs7fx0KN/zKClP9qDuU9oJxbfDuaWxQbn/QOJ2v64hgnnUf95m2UH/uz2b
KtPpXLHWkCxkFecONjiL3BH8Iqqk2UiWxI63i/dRI+0EBdccbURViFLnL+nS2p7J+fRROlECCLw2
78eiIMQhAmj9oLCuATrGZ99RbLuj82YGL56s4smroEkUmDZjN1KNhegu3fshK5l5rebtPjhiEBmh
l2cpkLvpLdwuxCNTxT2XQ6Szf8zMizIWOgWBdO2LwmGbd5SQI9CPJk41J00yPxo/iYlR95Ha1gw4
t9mlm3mmueUfR5Skl72upnrvcooEC+okKhjyDfXPmEF4811N+QDytMtrq9Xs/B9Qs7UfkIv7gmLO
ojimqS21Pd6DB+hgPBhlf3s4NEj97UJGoF2ZIYhcEkwK+2JvQuDUJgZ0+He+ItQytLFiNQ0d9MSu
H7AbBkOnC0qXpts9twjs1BCNaxEc/x5/FMGp5gxbBRyiWH9zJcZUYgCWBgTpozTTGDClW8Ty0Cqx
7U3qjEPsFRxzC8rE8AjluJK1YbW/KFT8oAk4C4gRdYBYHk8FEc7XkaRj7P1FF29nVfrSda4UHjPm
BSfqNWScSfiwrgZi1kjCVzHG92Wf9LOz9IuHFJKLtzX4YP/ZmegNc/uqzbG9QuSSojD0SLRTxBQ5
FKE3oYOaEUOaZJtbMMP6zd4YxpAsleCmA1HLozMbaJV+71RRFCyyjWM8Pj+3zi47MoCy0etuqac2
b/kiAwyHVrFIEIGiGbhyAwpmDjP0D/A0Mm27FUFQEn1vEgbR7n06Q96k4+3WmjlL2XQhnoQxBW7Q
lmM1dHSwcsPQUT/3jhmiLtcTegecSSSNldnoFnEpzt9LeK5FAQHlGp3AYyX8s5gQIMO1Dxc/I5nw
NuITaRHqMeVI6sDrWS/xSeSLRR7QXbZHjOXpDX5mfbQ6Fd1+hbWgZBESB2HGGponM8gjg3AZ7rSU
s3LiMYC49w50dqqzXN7Fc+5vOOzHq6MlbVGg410oU0h09AYdSQhESBb6yt7U+YxHfb5zqWOSejvp
Z1ZaPlq+iry3TiNftD9vLn0+SQj+sOGnSeXhwOFEWtUN57p/Wd/E1QW1WCjhIrfvbk1rEI2iKbZO
NQHk9pdMMbSPo5ao0fM1LIWZbMBYPtIKEyFaEwpesGLO0Kts5lzVJU+1GYTSnYM53/+yw/KvlAKY
YIsusZmploAwIMZo0cVzBgm/rAMzHnJwrfYVCSeq9+ysb6FmVef0/bB9NuGT5/g6FkXmGGevTTb3
DJFC6hH7kNazBxIPR6wDpQZVSC2fljm+pq23fyHgN1T/IQ31j1fdi78tQQ5SiS7KaSnk5bPQ+mK3
sVVGAVNYUAr3CpgpqkFw1jWragDHm/Sl66xQEybcm8eqaSVUZMEuLwV0wjb9u7KETeUWQCu2fZek
XChDj7SdToV5lybLTyvauC0RzQcDcp4b1s6T8TIKMf99cPP79TAAWmLXD5KfHDtvhEFVKSqIBpDK
PJqM0cCM3SAevAP+SZ+ELO22s92AFFIV02r44Ij5kJdasemjHGsEL5tpLscan/T9p+kj0bGt0Xfi
gE/mmtgX++RXzUsMyYWDKU6pnZYXh7ft9O5gwTMAbzP4KMyRBDghjeY0uQdk9pWozBcGEFM3hxO9
F1vQKdeKDq1AV/2ic60FQTW4RImwlY2jsZBXa2wU7irtyi5BXVLiQ9yGLaIXwvbe06YLCvPhk5Il
TCwWgYTnxZTnViwXf2pDiz3H6JDHLIAFZXu23hxHn5miusiWwmAh17KerJGMuLQEI+TumAPEilLb
kg3lpw6cUPSIMGjeKaxppI+Acbk9bK7mIUvNfq/gdqL+e90Iv7moCVuQVxdqtI5actDiRejE+gKT
jT4iXomOvGiqKMoao5myyFUJerztUjBLiaNOxT/wi+yyGQ4MkEz0aEPWBzRBCz+hRgapXHcE+qdX
ZcXs77lX4yg0Fo2eCW0qYMYppao/tF0ygqfQg5VHW9GfAb9Wps/yL3B1uvuQveVrQ10c2uVIJlf1
VOcpD8h02/JvkTBcREu0H6Yxyj6NNQdNzlvJjJ7Taad3/8l3/tvnWLi+HeX0S/bPYvI31C5jInmI
ezHglvCkSapnLresJwyZBk99M84GaRKk8PCPIu+UcEAeOeENWBQ6jSdC2nJ70LK73M7oab3Eu2Uw
Ng6vLhosRSyVu5MeDtW8s8ORSLvNTizS0GiHleV4z6RZI0vZErb3g/gBmk9i6DT6fTgVyoEvcUl9
QBMvAbva44nXBRSXP3PgV2VVIHh8j5L7pDXTcF2oJSIc4QGpMnd+jy/cx03u997yrhcjqXca1h4o
wzFz181y1/DUFq2Y00DMTvOxFyegpez+vVUtBwaAahmPhYnGLwvme9eRDeKRVsWTRAFxdkTiBhZz
BR8OrWZ4fYmZ9vYLEBS26CgUwkY2+qR9+hjBcpSC3QuMlMF5YYs1uaWXGf2dFyB3+zc7ZM1hYuFB
AwOtahQZ9uiapU+6AzJk+AWFKhgwCeyFKAEukF5os6GnLTe/lUQiGfWUPTRCPZJY5EXfP3bPGHAD
YGprzt4Ldzsi2g2ig18nZnt0VLeu4x4QAsXXoqE5zxNY/jFNYFnyxbdTEdrHOlsTJyBwIFKgmQa7
kY4UfAQytfp1cKujUp6esGj0TBW2l8ShKrflf4y7VfFidJ1/ERB2yryVhFCJQjJ1/PVxYMQk4Rsr
2XiKUELycpNOxzNPHHO0L6N0DyEkVXKZ7oeugZYF0tiqCagBfSTGDhLxtX4Ko6+Yr8v4nNWmqsIB
c+rPSyPQtbqHys++VNOIAN1YaF4T38murpdBEaq3qQi+u374JAbTFZXs1I7ZWhagW0m9qOaCwovt
IjGxWjy3FXzKJ6Hk51xFTztUvENEq6GMovQnhd3IUBaGUe5CL6eGtAZOCK/Ed+yjEcL5B/B3NXM8
Tt0n3OOK+ojh0CviX03OFaxFYU40ZNSsUWCzleO8gsHn/bFbIGgVoV2mlo9OOaPdkpkTjLkQwnNF
OD1nq1SqPf+ArzKK3dYm4ct+cgEtHO9piG3XhYpl7KzMCStvKF21M/TUbYGHjF+tbqZy3Rxg+NbN
jAdQK2AlUCRiiT3/A5gYPCSQnLmGcBHs0yHrmYzyVHYv+/FlPeWa2zP6dLQZuzMrNo2AGqH5sDWi
PaSTRklg0RuuxgUKINjFgIrphZsaK1gDycmGp4cTYN5RE2hVIAwpFu86+9sli8nmVCBgtNCT0a/k
8pNiAIdRij/KbpuRytYHs5XbzY22/Q5x90pSVv7+/k5tGZy23UytsFc+GDT8OK7tyCidwfpAN9yW
i/bAUeZ5mtcAd+JCEDOCPvAUKy5+GHVOU0phAIu5HVmX2T/ZCCCqBgm6hBbfYXZpCCcDDXzWvS1o
/Tvo6lgAg+TRsSXW+jBji1oaRAW4oZXvW5F3F8gJ5PHam5+m51LSuTFI8VSuucvQ/fJ9UaUO8v5l
30yGAko5UJA43ymFkV+cpsqu0cAvjvd5trxt78NxKEJeMHcEIJ1ATx4wkOolK/z7LpSK8T2AR961
0sGKCadEhgUodvqLuRfDD5Q7u++HY5GUuchH/HOwi+ym5vL9SgFymrLDDkH7cqlkzwfxf+hmsWUq
jQ+P09JpNdBIBmSzPIFf9yvHpa1xftN6UrXV0WwLjB2oq9dbQsA2Xe0lc4/lpRPGyup3v4Q7bJZQ
p0p28DOFbFap6SPCcgd1YDAJmKtaafl6jlQBqwDpMjf5SjF3fup0e7sr1DNFksfkAFzaRpWWO9OT
c1zIguH63inYnOtZdCv1ewWcb43ijc/A+hh/SzoF5ev1a7KRqYAHcoxECxQhgr5BFZBbqa0EtK4G
FrjIFhR3Qtq5DOMRpZgVHktVVN1tN0D7X37of3gM3w5QcMRHTxVR+b7JIf+jMdykg+/kdwtVhQ9n
2kIRcZe+fpfox5kAaMKzhU9Vvgd0N5LmcQwSsP3/l/TBLVw5YyAMOmKT4RAQXNgdJ2llkD58J/Fo
EobKEqeRifUid8Av76Z9kdtNGlMvF9WYQM7WJkIN5VSabRtfPadrw2f4oSameFMq5xRy47LaKZ1w
ZBLzXQB7q9NL7K18qnr1tnRju9oAKI6YW/bKAzaLnBME/QwFl6VddN9p05In18Ji7kaer30kTj7q
xbUgU5ZxwM9P7L9vbofwcBXiDo3wIOYojokAS8fW86JhPMkAtH3b7o7uQTvkgg15OgvxpfQBVAf/
efQXNHQi7FzK/BspNoGzbOATlOixkLSWxXJUW7xV8DtgBpq7yVfIxTd2Rwqh7h0/WGKJGOi92Wyd
Tih3IaLzs6KwlNT26LhyGy0ioq9POcu0YzIrVGvt73c812oouTI1TupPPlyyF6WSRib3RZLuo6tB
tTtuUU3OaleIk9uCPvZqCDsjO3PSdlHOmaLmUtQdmMMUmh7Y9dwDgZYg8345Wrkv3paQ+JGX+/gN
trumsptjWQ208qf3hmO1ReffzyDtxQ6AhG/z5gBd1byzZKnZJ0U38wHesd59xeMQeG97w9rJNefO
yFY7Ya8QdnxBJd5oi7xmJnNF9EtOWKBOqqjJ/U1CRESqfT81sK82lrI+z2hLkgL/aO0M7lTDT9MJ
LIZPmsvh1KQSm1TJ6POLWPrCDu+P4Pn+Rl1xhGn81Ca4W48g0cTDUYrnDKx3OeqmBVjJh/WmaML+
wVv8QWE86XjCWpBpSnJQVHl3Z3gX9FVo6eixm8gzATD4gFBTCXTtEczY8p/DUL6enR1RtZJG4bnx
ntjsbxsz3kVxs+g1ua3JGdlUvrfHWozaYAUuTLp+/S69NxA5tpEG4cv2BNW/Uom4B0h4FDGCqXbn
F5O/jQrlYRapytxz+EWENLmcbScmQiE3ofSzWo+ux6P0XH1TG0bLD0vZM2t82KL9n67TD69Cx1tS
jmjdy5xW+lt19KpmMAlfEyU4CHWXd8hCq+mPmLRZGYrNZKkIYk9W7bvg0HWi3y4ay+6RTFvvKDxP
yNnxXsSz4yccrSMMo/DsP7YA5DUrQdN6DCXZp0UEAOcP/jjO3jwL3O2cgequxvU2P7SL40Mj+hrn
olSHXtr42Jc9jOoKVUJx64ojoKV9LPkyI+Y7MWns6JBaQ8TUbz34oqCXpz4O3QMek54vENGqBEHd
nrj0HWLmqdw4prS76D4hvsfNTHsCo/nm8F/OT+FUvSgi08IazaStVZ1n8K7ANibDgGuSzaWacLAy
pa+kW5u8LJwp5hFnvnxMMZVj0WtXp6lS6VszzwfDtuDZSe0AgxY2q5RM1mhciDQjLXOY+TwuN33R
Q86xemgtL1rXbc/2Ny4fll73sDWsyKuTyjj+qLlfRh6EaAjjS2l4YiG8pOvNGHhSSFOliSdAjP4v
k1GuOPmEB88imckBko/BoT9IbO7uxNWe9lTLLMZS8VcdokXeoiVAf/19FBmBu1t7wlUeSQtVcSce
cPY951K0JWeYR4E6CUMBzmhSNFGEdOyLylIr8PR34BlKr54nPwRqd5oUjyAXf3pFCkYiF8KfD+b+
xhinLUYBkpfS14rvL1Enc3Qsj5UCFkfnq9zISwo5Sj2n0x0EBv8nhVX6K1rBANXIHaLbCs1FoHRn
0uZ6550crtcWoUf+lcGBDOAEz/6GXCM1d9FL2iRoIWQLNjgIblp3A2+0qrzaorChdCOiu+A9+j/U
6oKt7BQ07LJTwoIR5PO51f0c4tmi1dpqW7t3/4IOV6C8FTG9w6SwIWGTRyG8jTwIxEFZ6t+dBXC0
6Red5AfBhYYX/dKNcxpF+6IB/WemcU46smEs0ubS19fxgekSltUR/F8XVdHqH1hC9KNqQvZmECOF
wEQXI5J9yQ2kQDX+l/eUTljV9Yfj8EVBAWnfcy53Z2b7U4lTl+6KGVqk9SeUfZ45HiZf22J2R44g
QyFQ5UD1/pPk6ZxVMxNTO8EP9tImE1rNGHZ9qxrCYfm1Feae+It3f+N+wOV07fZN8zXiwo2IRiqy
1ljl0MXKFjZH4HdQIHpXAcz4RBHY+00CPRImmfVRN4OwxXSIP9hdddwalwP7lHZ9diLSpPNVoSVG
1QuqJW3iT5dQ2pJ+7sHBwnOO2fDiVl3FDJ1cMuu2itY2h1RQkS0J3MACbKahHSyYras5WtXHfq09
yum9+5FIndGpVuYFuNrVOJrYiS6NZm54UtemkBNw7FmAmC9ZqPOOjFSTVEPjm0Zo8rrbpheulFvP
2DSK+EN/Ut2CuvCPMHMrnwhwJSjhGjFhhAzDKYM+glumMSfBZQqrhdTRNXjG+VeL/sY7xY45PYfu
SASrfpIw/XtBwca0Ex+V7RR3Y/2TLqsH2LwUkOSwzkieM2Rfg73J19FLo9WGkws70O1m4teP9j0Q
ITYMkMn8Wixf8OrHwABXYSSyvy8ENm6rHmLyTNVAXrpsD8AzrS/2DXvrrNMf0UVzLv035wqrFMl0
BZi4Cmg8nnL4hDFpdAtOAG9LLU7FiEkXIca0yT04//0JDx2NH5O4+9GhiKGTSMDVuNLbvXIwQ9o1
y3OHY9ndO3pE+ZCHTNIgiLzjIXIF1EUCM67hhXbuVWXooGSbQVkQfRpMxts2jcj6O6DbsQbl5jBy
tNH+TW+8Wrgt/kKZF9z2OKN2KfnXyQ/r0sGbQz/K2Pqfa0Gjs+9JK4W3FYEbL/bchHPbd4RNKWMP
XAHvqlZuci2qiGX6Wmn0nZCFeV5sEELAEu2oF2x2NHcc+E2ix1PO0I+YR3CbwpK2cH6yK1nzdrRb
zkzNOLcaTpaIMZDJH0GOs5Kg/HqYsGUhdRT2w6GR6Ac1DoBHGPjW0/15VDZ+/td4II0CUT4ZOmUq
8xScUjGicJTLD6VSRRpq32tlxf6gISl7whAW57uMzleWTn/dhuXxUPRF6r+IcyD+7aY5UYBePV1P
Q9nK/jrJa2SWrYVy37fyuZr1JW2/V+SglAVSi36MkUdgQnnpU1IFlvVKoLs+ubLzivYb+IztOupg
W0/tr/4BshoPH9V/5tiKIL8yEE3MvcsWovGhcimVZdmei8hyL6buB4KUq08a2IeTW/FtWzv3rN+3
NCG2NfItX3nFc4qvTJa7FNcb/StZb5yTl/FjJ/HhWGX7GkSzi0iuzgniPoop7je/QNPuILz90Vc1
5TpPP2LFutEmRfg4legl7j46zqw+TBAvMiKkCN4+wNoxGXVlA8XAgqUIM+2fZhlSOkwcXeq+Zaim
mDHne7/8KY7KQqsiHdouE3AXfUHh3NAf0o8fMjmXj8irSdkQf5eRSaoL/v4/SEvLB6pNs3Nfiy7o
AA3swT+NlBYhb6kpnfLr1B+plcDznBYBMCho3taYoT5nnSwAWu5pvsIOpP+Vw4B4asGhq2t8T95q
EzRk1+pYdrAA4YuYxlO/B9DGzJExRpOpeLa/O+vb0T3P4v8t0u67jUIMCKcMIzS4PaSiYNm0RFMU
4BDL2TvjRUmb/n6AJRWDwnXz9RttfyaXside846SG7vMvGmoEcMjA9V8+SB8gA5jy7eagpyH9kE2
cHhbTC/A6SJyIIMPjetb9zzOzuyMr6aW0PMgrprVjvLYeCjAvQRc5sg0t2nc1zFJuHv9DdiyMAXG
Y859yiW2Bpc18P+VgF3spp4LC2oQefjO1ehPk8j8v0Ici5mnUxTL5CoryAXKHQFA8ujpCb1ooUPN
YRWT8LqafDRqndUh/+j05sRzc0ZsCPDAyxNdx3zOX6YklAE/eSF7/+tg/FJ5iwaAijCf8fQPRlCV
Uo8yokRGjpN3lLxdxyvtCLWxn6fr/6tFhE95swfbXrv6kTulpyRjUZVvtM6mCBC/vGUFie/lH7OY
aYSW24tOvS0GkFnf1X8lEFjbyp0kYOsTDCZsiKY9PHt+GzzIX4oJoJF0prwNaR9zHJ31FtqcR3oz
heyMp7tAMeHUg8YK2cV5CF6P7gJxnXUhlMIxXE+u4iBn7nZUs/BiBSycbmBnoyhuJFQuo8r925Vw
FzLgdXnhdbNUMBUDZVlBGb1wCneWiReC26qH41SgxlfRqzTpgjKUrwSkQeBgzZPvr/x6gYyzVmwD
H881L9hzm4JqAqR+fD8Wy2VxDOijKGNrOlPuJ6L+Bfh/5osGnIzZPic3tC+lxR4mepCyZbeVn4DG
BxnqZTOtXu3WOx4uztRPr4yZ2c8OQeGyEAOgKiLIfHENEzHWn/UK7g7wIE9J4MJSs68yY3Wr/nSZ
Z4RUUOrTZrk0Le1y2FGfUtP2oLMytPqZmbDjJ6DSo9b1nY+PYHxuEgwrAEUmbz0d5NAS2sXjqBr9
ICH3AUkUe1C+SqgDycZXxhK7RL6vIgFuPgh+fZWTq+b2+p7kiDySkDPyga75IpVG2RK4akcc9o9p
97OULpRgSmJgetJZ42rmzR7PV3iUTJ/HV/6k6w4SLWm859X6ep0l3pOIjEB6a+gYsJiuZhXwL+yW
oTgfoZA28sR14KtmX1ZV5FvbeotoLkR09Yh7Zrwtp/Vp0rumDYzHCVCKgg2A1tqVBla+hYtTheiw
Nq20cd5Rv7nMc0SoPl3T8fYFS7nwaUGQrADbAYgwqxDeINrsIALvj3vQgtvWj8WD+2hUyAlZo+BI
y/HVADfdNgFpGEzARRp7hYs97ZvL0vgwaXS2seAbhJC5Ygt6A4x+IqE9k3oslcwD6chsRgCe5gAk
SMbX08BhBcX6d7Y2mv/ovFOT0Fo5+m9AqHJnpnFDFbNSn2tnICYaNXWbBwG3nKQXGNqygdP3ZcEn
9OSVfzNPK7qP5Yzp7JOMqLcSHsu+wk6Gr0FKUNE3XWndQ3YtZAgWqdrfOUWj4WONAJ36oXvFe6Qw
H4JdNTvBLF8GULwq2i0TL/Nwam/b/D6Kp/WOoex4y7YrPXGB7F1iB/oN8flcoKdFsKquuM2wkRf2
qqZoacH872taFMFSSvxVtImezcFlCC1qUt2asE1O05A+hr+5I24OowiNFn6goM0gArRpqlUKK5e4
yPNOGatVhlRF2m8XB0qmb8sN1Bfl9GRtI+5iKn2btb2XXrcCGhANqg4dQI7Whn5E+9wm/mLjLf19
rOJL8FMITACBXV4/hbrsMFuVABKezNzt3URR2A7ORvjpGFMH7kRkWmnbatUeMEi7kOdG93etOvOa
qpzG2Jywa7hHChThrI7jg7VWeVYP4uHUjl0FnpU9WOM7Plc9qFJlB7p06fgmbgTFwNgY09e57CPj
r2rMb+kY1QUq+G1Ft9CDCjFgLNSpTKQ+3gm869859LUzpbLa62ZxiAzfF74ThUfhPaIxAbJ+6uyI
LoSwEI7wSYvt1DBV7WoUMh5UfvN8iUP2E/9dY19Ef11hqpRIfhY5dXQMX4EHwsX0u9ZAc8Kshku3
Rz5hc2jxX+wbMiufNdi538GvOEpYKOGG615tD3J1l6vN2IFQVh8+vMRN8RbM/EpucrNzQ5tG1ek+
lC4HTUYS8PwKKEF14mBoPTW7CLZwocufXBat65+v7jUuXLu1g/1Sf6D4G0i1SEmYluk55OP01F2/
v09KFSnShyFa3xU7t2IZY0CUcnyYr+S5xZHspYz2QLhg8nKjpgdvzxKFJaGmb4QPqVhvGU2R4bPK
T+p7RKqnQJ3aOv7gHx0oQ5dlo+XpZTN5K+ND7tLC6JLAQtd1MI5ljWkowavzoPmGSQK53nQ1DJEu
M/CQUqe5Mn4Q/8gZhQdwLK9AJ4FnZUGp0TNoC7nJVgbpb4ypw/tE/xNh/7DRts8W+W0pG5+9EbHi
JccZHJBaqpjJrdUUHR2UgKJwhI6+5HPXehshDETslSje5MRS3qTFYqCPoiXG64PVQ8rJ0vptplKb
uUONWDZXFip+VEGB4PmJUk1/SohIBErh58iqi35WZOO39HNy67HnZOmdncDq6Z88Qdms2IW6nLYd
SWxKMR3udenJ5J/zJfaKGDDfPWZA2UuObcb5Qt0oD9n8RCtrBh/6lCVzFK+fyHm1R627UAuC6VpO
GhzmHFtrOfA3XItwkc6/skY9RX+8QQnjUX6NoVQN8KMgj6+o8AasK1fGHhA7R7cQmw6B93vTdQsy
pFtl8yM9PGsgNVJqkg2rBlkyv9nvc6nLONudJBK26g2DLcuHfu+9z1kE5P/lMEM50WD+/CspDrzr
AgQEyfZA7e96ZLiRI847nw83Oox7rNCkGk1s5o04v8i9MTGW6U9ST7nk1OpixofdduIrbWs/uJCj
4UQpsV0zYy2wZvBb/Q3GufSSEofJtAN9PZSVkpZogHXd4pdIiKY+NaMWrsahFZ3sQPzvJnfFCtaC
Z1eo9k5Jpu9yog/Vq6HWn2gL6dc0ignSwthYBLJ3cfUKFwz+uhMQs++xAAfszvszKmzcl3hUzqb4
HhkXAMa654JuCuvthhGnLNG3XSmqEws3ND8KB5C7PSTdCTWEag5lMvQsa/264s/ob1J0Ty9IEAie
sJzT3ltoXhdaRR42TfIViOzPUOJeTy9+QaXFJhLxjCTxmAuhRUeohFXwGW2Gtxq9WAA21nSdU7Z2
n/GqqdZC/zQGEy7GLcASE+9D8wLWDq784Xw1oysMy+JVOT9K7thaIhpJ0l5kM87p09p3a6LNbhHk
rV3IvU8bErV6yv44FA7YhlqZv+nCm0F1FMEbSO6yJSCS8Zl5sgoqJq6UWpNBpkRQe3Q+tZ2PU6oi
P0U9QRtsoJTr31FQyztUQkapQT63cDVFUn3L5ulJ6lF9sIPKTaZZLqsAP151OFwxDEr/eun8Hk74
HaLwMY2e3hyo8Gzibfs2gzzArNKvnrKAjkADWBFs4IXZCs9UmguvUJpGG2XNnwOgBSzzntEvNpbh
R8Wl2UsDP6yFjsKNORlu1kXgyzrJoJ0oipV+NappBZTSZN28QusaBFVlCcFiC7FZ5LuMAloNlojT
KvOHKyljE6Pg/vP02BGvdVxdzaV5kNEFrULA8yrpf2gF/r9Kl0KprBw3BwXLM0et3zhUlYFh/wcZ
HReZUSv1mz53/Zh0fyB/X6NoQLyCZldfYss2MRChrCgalCfSEvJ41c4YzuSZ3Y3R4nP4Mzsr0qBO
Ulba8yc6nJ1RMZ9Zvq2KdzBxOTUH9wRnZYtMvRzEtqzoOws9hD+3u03VOr5oB4ZF7CXoFVYxIlB3
dPYA2GQn8imsoTtOqt2CYE4fEd4+Rp4fa5a5Kvfw96efevp4Aimx3/qgmQkgrUS3dS06px/JdajP
sgMc5evc8jMC38UbwdLMP51nunegPZresbpNdKa6QSPa9P3PGShiQAd9aoJ/mTZ54XBEhtvKPn8a
n/OcuTkNJQPB3lv5ehNhU67XAPS3P5W7+vGz7n740dHJ2rolgT5KApayEwUt5edKjEHXVYo2wD66
EdAhocC5F+QnQnIihtKP15NQRh6VvZt8DD5QjAkOvP6IVd0CxCBr4hAT0i+rj7fyZpM86QzySd0c
ejuque44k47nT5OuwdARhveZx2yWXWcqLUyC0AVYjykOzlvT/jDimYcckojgR4rIQqDJJNbBB9MZ
SZKBrM9dwYNUkB+Pj/gNkVgTbnqr9zWoOe2itp3F8zf0N12vumvUWEiWdVRQZPSVgLvDBcKJDlpe
+17gO1Hr2ZyE1h2wzoJSdLWq9ZRGr/UNI4iBzLb/rxT51LetK6P53rCbrQ9XfCzUsBCtUHBR2dJW
91dWZnE4mP0YCoS38SouRNxCjTWVvyzSMv3W3ZWP3FOIBb+2TD2JyY+EreYp825Mf0LR/yu1Y3gs
+PLzN8+pPk9ynlrqv+aXER7O9dcK6KUNT12EtIWtkbOk/26P3NMOrd/Z7w4T0di/lsCIAS/fjZen
1+753FODsByAk8AM2Adl49ZLDepBL/5eYFWQdH5K7IXUZX24/wq9nYbYAxxETAHN0w/xF8XUSxYs
ZVK1K18UpNaxrqHsYVQ7sS9dnEaQ1KCss6hvSHnVgCPNsvSdviKbRih9ffO2hNu0yP3ixqVkylX4
NzelsWzzrgTLukTqgM+wwmsM2M2jqOiRXYqd7yKOeWQV6jcguM2IICwohm6ANgGGAvhyhxloPZh1
AyrjFtdQ11QsZO6cE4us6Xkq43CwOAhsVGAQ8I2iGkc3d2uU3OG0QLawBxWFJOgMB04VC80RJ/Jb
xc0jDSAF3Jrs64ebUanbMhSzZvaaVyyMzcpd2glADV64ikCjeRUxoxOqsTyXJKJl0ztLFql0ZOY9
yijnIVrPUVJSLRimSDXAB22mDrKVN+oXxNKyWa8wgiBJqRRnN6Eb9UAi/Rq1qjTLmDzA9rggrzO4
RyLwGfOXjkYBFWbXBQj5CQgvH9XNYJkI9wH00pGUs8LlWikk6z0imY2owwlIu3Txt/SofFotqRFn
vMoKZGg88aLfez6OMGb0M1f3pfa5AOxxIuhvA4GHSgIbE1yYxMbLV/hZQd7zjMxVesG5i2szLbx3
Sh9xMCxVdSoJll91kL5MbcpqzYdknvGiAYK/xXOX3CDRGYycx6cZrq1lD2rcgyF+lJm62kmSm0wA
ByPzWa10aoC2QHizdyBHrjqtRRgQz+j1fm1bnxnpgQ5DhrNlDizFWPvblRFeASxJTvMjQH69BJLt
pnyQekSxRQQEKGWxNUvbLxd4K0hU6F6LTXXGGGHNk7/Yvanea4pXNVftlC56C1ClkioW/9n4ERuH
mBVOd+d++BaNPEdhopW3hymri2Hpf426AScmM0H4fq+ytMal7T8a+C6V+onX/c/9M1auiJHIgFz6
iPLQZ1w6MFYRxyHX9LNc255AoaK01NtVHvkUmsuTC9EqoZguDMJKWdtXUnVaaGNPqpX55gE1yOL8
wHWwKv83fpyFbhq2o81WHoxnlqE5ctXiZsIKkeKyo0E2/RJipQnb3YMkEv1BOdfNsIJM0QaV6VcJ
ggBzl2/wZky7mwDsb8byMdOa+FC9Lco3388wl2c+zu4vTbq49WFKxxdk4BxijBw40BiEOcMVF9Ek
3IQZKXfx5Vfq5j/oX6Ze0KcBFR3Z7iiTivGAnQIFlm9Qj3CiOzob6e2tQ8S9g61ANcZIwHQUeeO3
P5i8q4aBZZE5/gwcq+p77VLObeazgEVPyngExqElV2RMrujT9N4arEHigP6rvClib5sUsGttTKTL
dYVSnqPZOxFzWUsRqkUFHVSlJ5VxQasY5CtJL+DPLkScvVVVgVHYLBWBm3XC3GSOp7abpLYDLxhr
ZG+Z9r04hgiC/rbz5kN94uCBCYw2b1/OB7VVOna/iKS/3Z4ombQ0IeJTfwivTzbCbyv+jzuq4wmt
8Qk+yS9hRPqPU/Dti2QLTqn8p+GUs9E7zZnP3e7HsUFYOHC5HDVaOUJp86iYeXX1sUmYCZ5cjs4G
dpEWjIe2UzrAC/Njl7Zry/TS8hBj+MABPbcqHc1qED9ikKeikUyf2rHca2yVPOOqVCIPdtl9/Eyg
L+b0UkX+1Fkq2TEBFfDXw49ky1FgjEI6VWLL1j9xMf1gyP9hz9PsWD4q4uRE6xQpTxkQEPaMd4Dr
OW+BP8GZD0itdUbJK07ZL2fFIOY4mmed0EzizVUaJplGuUjz+Iph5oLw64S7H2/63VQI9aUZF1Cr
9ElI36PTU+sKbrq8jaTp+HR+Zn3ujP2VwGKbVfe5kSmIf5ocWNlGoeA1zCkU4yIvzegYQqQMK4/O
+ZiDll/cWVhQ493rrKW3JfzCLRQa5mFd/0/4RZ5Wl1Z5sxYbbCPfrykoXVyYi0fyt3xWaFBLvqvv
EgN49p+bcBoh3K5gqjFEaKR4Kj4dj7Jn2J4zDTh0yKJjBcvLUjp9pSFUTPz3y906ntgGhLnL7M+P
vT1UUgiRyRJgGyQ1QXNTJr0QK+FL/h24FokQMRtHjctBAggnI/A8xvPUdw3G7KzLV7dOugqWg7TU
Iog3PFZqeWBSZGunpCnMl+dxkM3wUdolhoPqN7UBHAfU8PVZN3Gxb1nafnTqXdOu9sxR/mZgexVZ
YJpZbWvL0dz8Ns9/Zqz9FMfm/jpFO6XXs+5cqdDocdpT6Zppt9iuoeDsqSauiuMuHfnwhxNQRzX/
8os/ufRQDw3QQw/+6sSB94ZNHQ1qB/kyCRMqeVT90rsywRVK9apiF2oHh47qANTyLJcH4RNwpjq4
sBB+ZreVMKKlqP+MbxfjGsFmHGEJ6R/YydxPXJoJTrQ7R3K8k0Qt4NDlaU1h1/CJSUMIdRGZi/LT
aiR1RIGLvmtDetCQSN6zAAa3X7skodKpAFaj1wi2fEqcdKGxFvihhgR4cn8UuWEvb3W+/Hs2W1PJ
npMNSIIn7hmGsOgvyxEP2qHCkAYYdiMKsd7qAWCeWuoExRZAD+swv5m4UNjBVup3dMrm4QrEEGA0
voa2b0ZqXj8tGObzX/HCPPiJY9wMoLcU3M5fs9L1mJpx3YgK430YlF0i2rogK8UyMKwOrrLS/dlR
ezdbPlvlHFhR6P2UgDBJlMour4v9e9zOtRSUDCM/8Gq8kL+JdJ/DvONYgqBOWXqAurgLbw6JMU9I
4JqUT2b8MptYCKeKJ3NUVptsrHqmGzQvUxH8VqLk/hRCTAc336Z4c3/RCsupwrhYKyvLssZ18p/e
vi6jCTNmOiavUET54eqHrGVruTfpGnJScZkaQMMhJGTlh/WeFaFZg5GMltEeUoEvS4vxixQ48Wnv
uEgcCReU8IRIr8qv8jGfz8qu5hRGBOg2KzDRuNov80Dpn1QBEGFyfutFdLYjw5rfmR+hZHeAfYv+
7RDnGUYHORe8JDHcnOBWXIOFAZArvt0gaPG25bpFmbR1XQVODqmCtH+Ay3awQPF4VqndndH+XGQs
b+Tjcx+CCBjMKYfLu1k0ywwbokRJ5rfK1CDtktxYdXtsvjaatq2iNVVQ4H57/iZci7ewSYiR77nE
hcRpaWfrdxT6/8K+BQlm/dtKuL7Flihy3uPqf58t8UY9KP/xrQoyc73UhVbnQtRteLHoGTCQc2TL
MEDK/NEFQ7NXkq7g6J7EfWkNM6k5iRfS6aYpHOuzq1LDF73iWWSds5e1jHrZdOX8TTIaqdLVN+el
DTtRyRgV39IwN+OZd8y5IgFRhSfRzqYuJDV85VS/taqotpsxHU8PqmmclqjLcM30xXQ3kd7QRhCP
0ixnzIK9G45EgPyELMXgiqiUngY8mZ1asF7NqGkRe4XSAQxU9CdEwNpoinJDvWhHNCZ5aWpU76Ha
+4xSkDeZNaoWoG0+HZe8nznfi42AkDUBTegjzrhoTpx5llnY7ZjFhGfTzf1dLMkNK2DaAuU85WS3
PABAfydUu4Ovl2JuwZ2FqvXpPjwvunh0329Glxly2FhIXw0oxLKygVYr4Zq4MwO490JaYVRDZVnv
s8+lu3MWnloy/RvhiUDEppwACFpT1sm6X2fay92oKPvziYuzC7IMoBOULutcW/4Q1ln39Bb/OvHP
HL0KjOdIdSodmp4mrdf/8L3oBlGvY/rKZ4oaYZuypS9IBceADrOs/h/x8igpLu5Y2KU8Fodscxym
jXZYGXD7sPHRIYZmgEkeLzA1dohFwgFmu8T9zADSm34dYqV+1M9gVxyrT5gvBjTgLgw3Jpg5QWQi
5FiE3rm6hWvXr3SUWV7c+DQCRcoIwPfXEKYphQU1QA/cW7XcvJ8v7LGv1VaqVEm7SmTCi0CuKfbf
lCK8y/sxW/K9OPgEvTM1vWmYJeNBG7Wuzq8JVwrj8EwydgJFuF46690RJ3SdVLJVE0Ip+m3gsyXO
8MV5se3/bSoqSL2QeKHx+FbOJGaaY2lffHZK/JO0FZAr4IB/pj4+YzMgzmcX3eTgooZAh6HWutHb
6G+rraz1ALCeu79rQ5YEOXcgqbsp0l/7dy2HqIb0mrPAB10vk2R1IgaM50Bbpg+HfHY+NGnIzQxp
oRWfdvY8izE5H3ojQL15UvYYBmXPfind1HVCRtxx4enZMWx8JNjDMh5o4A/MlZv+KRadTedV7XlZ
6CwkL2evd7GZLG4A34MW5J/z5DUdFC2c5rNX5I05/es0bCc1sKPHc8X8IdwLiTt8glCOGO/uLP4J
Cmg0LGWcd/ji/tj/tES1HeNoIiE5/neZL83xFlCfOpH/sJLj3wX75nQg+CHMelNeRV6TtloekpLa
eFUycDgNtHtXrgUmeXrroUNqLPYQ7kUFhk8wu6BKeIEfSSx1LJ76YMaJQCliElPRjKPyij/vbXuW
B0pNE/JGt3OAHESMruUbxd/DkJHvzOQABwrMps6axUL2K+SO5HCQt56MjBMN9iOckU+l+fsDK/P6
SxwiRQZdAXKESl4mKS4mB5pehN5CFs8cfIMxJHJgp98nZQkbyy/XF6GC7paILeI4IE4krwz+BIQz
D/gMbJPVakLaJ0h1ok+ed+XHKwHJyoyAStXP8kxah9GMGVmH84udUl7OTU4AWis9MrOJhRGy0lVm
KQ6mcx2SYgIaKcKMat1/qAsuy+b/O8K/tjEdHN6TtRVNqfvLf8d8Q7mOxg9uefJwKUCdvuA/deoR
6akUvaux9pstX1vm0ZfJouPPGhXpi1e2MVes6a+Ld4TV8hwXdCW8zxb5sBEEp/fft8XDp8LXjpxL
zNsceamR4a0qKGY9AjgnM+yxks6n6IDVg6rxHDvHEYtedz4qrvwO1lHOKHO7DyA9ImYn8H3BYQHC
JpFgLem9uRmAyeaYGR67CA6UpyjDwyzjvBEOYkC6Gx42OrfeNjz1mXspKFN7JgXFUlk+ixiG5xps
PywoMCcnmb7AczwQjlv52Tyu8xEdcZ9UB34DnwXXsFYQj1OXSGMuX2XNx343ABlWEte8L5HpKasL
wfEY9gk5LFJrwPbEF4gXv6+u3U5eMVPJrWNEm8xem/oarLGry4gLHqSd322rzGNWlD9szhEHXtSv
1AuwMM8M4aocS0bPFGVjou4MroF2d3aErmptFrOKP1PXPIFGFNQ+Yyz3DT4KnW4G1usxItR+iyNs
P/NbZ68+lp7C913Co5OejycCyUfvGYi2p5cxSrm0uoIo+gNDn4ZhtqAwOt9KD3+gUrnB+Pkl3CqD
6jboMXSidfL0c3S9gWY2Lt3sLECgLG8TL4lJ1SeePFQy0Au+87KWZ/ZFLlzYEvwAxgmUD9fMC3Pt
QT7fKtDLJ/LWk2mfve5ntfELmVmVlDxU4APQW4dRzMSYhWzRdis/C6KZpJIsXWv6YENg1D+5btDT
nhvWSognc0CSiDJ9jkj0YuqbE/X7Zge4/WYVdvQS1dKbUuDmvI7xrA0oTQ/sH+GkDSOsTJ1mkwzr
IBz8dHS0a6G/LLjF9ifLhi5lhcvnrm7nigZrQtlPYnPTfyIn2gPkmE/7mQ7eqSDAgbMYj0wjXVI/
kHavoazzB3Z7eP6Z5UCUDD7Ag5H1yCTXgwH96u7+TrSq58nxBhQNB3bw8uqsgI22UFHby+JpnZvG
NtfVXXpkGD2AxqsUNrbazg1yXH2Yb4nLmavbAACrWJef2I3n6X58wwkokyrMe0VqBpGZO6MW5Gpb
vsaYKhG0iKI1Qtrby3P8wNjtENnumXFU55I4emSppoaHH7ClcDh2MaPTss+ukNlxh93vSa3CUdmf
EtafcvYBJDucKLS/4QIuxDK6Oy0x8qwiQUuUKklTGWour2Z7Cm14e/mZEUykd//TGSoObpve/GXO
+pbzyamkAARXE5anUzjcMn8D0GYHPyTukj8yVntObT3+3QajP9qOn6ib6prSXZK40pLKhIfvkWKl
IGXcwfuwSQUH2b9PIoJiFJSX4tvS9g0x3p9SzmI9w4pEmlVISJ4jgGNHMpbBWlXJbH5axYrpKKS7
FK6nYknDAal9DC3IbU9Gj1Jqckrp+xf0O0rmlQVTQpj2ijEegfeb9RyBPR2DG4ktFv9uQiCFors4
89qHDuv40Dgrhxd0A86Cd63pcCqp0yfaVatyq0tdW/672aKb1yj8B2JyAN4etvJ8A5bOMvDf+XrO
MJNnfY7lBZAq6HD55PX0Vym/q94+nRJ+qyXEYrC/8mwp4KP6xwRTPrRuWS7ivnU9vRlhWkAJGKb1
jlv8WLi2pCMNYK1GsTKlm+Pa35rhbJ3Ul1gFNyY+IJNlqzc/Yw1qTcXv0kJ3QKUWCrxDB3hZe3mN
0ZEJMeIY4wHffUUUr1o5L1a0E/jnCYemCUwou+sbXOpNw7MTZQIIDhzOC9docd3BcHefRDmRT7uE
68a1YoG23f/UNPATadQ2l51Gw+60WdD1JbxRG4OFfC1ZeJeYSBEXE3wxejVvFaUZKKPseVY++9O3
5mLvd+R6gSKnYHSr1TIK7Md8zhWjvfVTMroAM3ax8QyJgqCzwMVNaBAiU9hdMiUNTcFzPllOB9CL
E92hMM4XGXAfO+0xffxHo/+2uU4v/Zkk6F71eKevRoaSjZ+joaYqHa2db6Oe9ZjPigydlr+q1pm3
TTvHEk3htloo2uU++cCS/9KUQurEoxTnwyXY7t1gWFFtFWVyszDTpSxaFtxt2cfW0VGNfHNTqw1A
R52575g8aRjSKhMiyVhUTS0PLTcPVbP3TFFQ/HwVs4DNGLU1NMwYrAJdGYf/if6H7CW7D00yktyJ
zvQvjaEFMROIWoqx9P6GZOMRGYklqgn0WJ0PVX/w2NrVt6H7QTQUnu5ZfqluO3r0LpgQ2hFe6EP+
7z5WHPIlUr83tZw6NEsQmzus0Lvj+mTASCnrEF/LSEKch0cd+YrtNwB+g0fxSt6wYFONsrsFkBaX
tlCLINEmBOycA5AAZfz4Ng3RNueacnQ3AUVvmKCBh7Ye9c2A98FBj3S5taVlDJNqho7ylqJxQ+Y8
BKh8zDLYDYY9mgDj7Qda91waP3lsbmCnSDRKXER/p7o+avgXQ1zZbO55qr53lxbj2aTXQ//Shnpy
BIWMAAjc4H5O+Mb7ce0lTk+m+pYjLWpHi28yqcuuXuV+QY/uNWLCuec+/iRTqb0h6fDdT+kD6yLR
jBWaJsHkQZIErEiqwJ0HOXiwNW7HjXcJjLh+y7vR3esCsllfUgaenkX/t0Drvb76ADyZ54on9Sau
1nw+yfqAE7G+DRSQ8Gm49CXv9oiotybCPCKgoZt0bc2xZ/P1XjkQ886D8jQJif37eatJNZihgzhW
EMRDeMYirQf879Z2qBKW8PJy9i1BNQMJ883fQFTdNOAs4F1oCTHusaaB9xu3hhy8QZmIMMShQIGn
0ZG0l2fF2FaNZ0nhCbN4TWGPkWYSNzSPOUVIkK/u9vgSk44lYlHeDFuRh1YFNtL2dzh5Mw1uqxpR
9QdH8K3+9IMTVc06hfHcHmCiplrLAnzs+kUImKxEKqJ6VnDjNQtoBhA/c6PW0zVVuxZ0uG1erw6k
dlSo3ccE844vrgimZ1dKBOvHUoSnQ2CdTKarQks46Wv+vboeKRqIiGtf+H6DHawgkWlmRewOGhMN
A9uN8WT9dAXHfzTHfXOjzsuD/jvGtFAW8revWTIFU4HOqF8j+4tYLG/MiL4ypLuK7bCraK+98KdJ
X+GI0O4Q/eeVQriojed5AqcwHm5xXSinZvUyW0KDfHwhc7nCPBMYPaYdfwlhVDkoQS+n+1jBxbWq
EcdUhzp1U8ZUBT47fl+BG6zbmd2ZK1xxX1UEN5EOvJT7VqY/3vFPjGFx8OZu4ywOg7XDnJjx42Sc
DQheFsbTZ4vAhcQPNj+uweW/uCBKYxEUxxnlNxKCS/16AJktTT+7u+KxgGLR8N0CIidBTM9auOu0
i1SjRHEZk75QUZZvYRKUk/tlr2l7JlkyOpnO1TLTV3Ey5q6ue9y80G6s/ZGrSNVnGWEz1WDLBwxc
lVADOyZGlbtMN+Pj/x+DJlwOFl/9cSdQKMB1tOxE6gy5RbrX01aQ4ojIhTVOevbdGjfuXQzCsG26
Cy04LK0CbdQV4jdeWVrfdPpSB0wKmGVEo7vWutN7GX837E4JMXlj0DkMsWb4sFJWJ4MhE68eb0zX
qztXZSNcz1E6YUmJhbUpV9f08Ornr3Zr9gA8PCh+5yDCITA6iE5PUXITOtsZky1lZew7MZjtbWpW
fWGJ9H6lO6/lv12ACT8BTdbTvmcmf+5UiDf1LZBq4G+neVe9KDXOAmbLyT4EjXukzshJx8eyX1KG
tT+K1yqvYQfQzOkHVyiR5JgKarzd7CM3qeCUbS3NjjMhnyk0M0HfW1MJmdQ4HFWLG0wm+3CmihA8
rPdSwxmoyvNJB++yzk76RdTqEwdsd1B5+oi2w+WGUzKvrjiZqhsg3iNRMjKrl9GUwVTbmIdoh+M8
4zZSTQik+zlrvw8ZcCzGlBAFjP/rvu7HGLtyJFSMCxiXfEzNeM+gLB4tCV9brf1xaSnzmGA9ZnKZ
nR2Akf3jqRJEwT/QOntMiJIXn4CxLdB9+CAPHsrvPcRVtWI1PQ2+UAOYxkuGV6Cg37vuxF6F4TEw
0Yd9fl+6QHNFYTg6pWJMkPsNNr7gwQdXWgnRQiJzXE6JJbBqL10DylfKZ2xmWwGa0geyDL77AQ4H
qqH1zDIFWUOiReR47ouANfZUSOx2Al8zpTgy4OsSmaCWg6gAC/Od872oCemos+V+QQ8xXsp6EUHL
AIswSy4NN2M2FaCmTCTXXlWmVOYVS8cOPM1CEafBU+gTz/JJDIk2L6555ZsHdmDKnh5a4ezsSmZF
VBhzbaDPb/lykwZg2F92LQTLKub2AYvUz7GqM/4J6AOx+GTWwFrZzIfZjCHzZDfrXnJ16NUCCbiq
+zEh6tHGQWB2wX6ltCgYjYOwQJyUOxVJhQq6R/uSCZ/1GUPAu8LpNaI1FJhPvt/EkrEHEvC9a8lp
Z/qWGJGfsPbxAcz4gb0R1SNNjxSupm4wOuCY+ZrB2OhyWXkAoExg7mIG2vjxoh99xsddxS0G2fRv
GNDxiMSNNErQGx+1FHTrpr7AhYjEHTaM1BpZGRUPHrEaEylkDDvsan3yzJe0AquXcTBy+fVHSFUk
S+cy29hItwTyGUCkuByCbMWlWH02k9vc/twefR+YxuXKuTySoUfUBBPhaOAOO2CXlV2966Owf61g
+t51QvDjeMT+EV5AWYobGLWG0cJMmh23yg+K0wNP9QlllhFkdcRRbMom+q0g/ZYlQXelQjftJ1Yy
G6nsnGh3ZvZa51yVRJIXjnghuzPiFxvdgAKbxzX98YUixov6P9VpLH2Xs9IDz4usX+ZrSsHAUAJs
yskRIPWZeHvobjDOjl9wnz+RWDSzyx1gXCYjHibCPv+khgNEAOTcLK+IxuqnI80mbfG0O63oq9V5
i/WzDmEqzuHo+zvfbAvpRVUIAN26joayGyM7EeHHU6RvA5fXSWG9QEMefe4WzN6KxXXNvTrtW/zw
xU5WKgCqSnLlIBN6BsNGZG6tr736OcA1HcFhOCxgjKBMUlWoe3TwOmtYacCi+IK0aHuuvQtqIB7n
p+EkSBw2XNxCLMfru8bebgQEA5wwA9eCubJcKN+pv5kx0uGrczJdtx87gE7b59BTHRPqTwvQF0h4
dhaa6vnsaKIwPAkq8RQqkHNJ58KC4dJpK6dDweDYehzEY4IYgnwj63OSPeWuff25FZ2XOKRjBQ5y
KSxV6wdDr388VnKLqWow7EMFwATkFQX0dxFte1H0soJ0ixO1OWhSQoVTmYJ13Tqn+EpAEmaDGrPf
YKazc9cmYNomOmV0XJCZ3uxcsP+/ZoBuCToskjcSXpjSyU+tBfwRngaMvdEq/fHYaOjk6URpuh4D
NeEtgCUVnPpNk35r9CLT0iHys/ZPEpRVNXx++uBbUh+4IlMutQnuRHKaWQ7ZGPum7V4oiO9n2+7n
u8mjxwIKNE7GjLUYzgp7+X142o4l1TtrGNUq1YTMp3Jie6wI6lSfW7QD9BKUuDxliLNAp5t7RTj/
3edT7knYwbuxoJDFHWexLanIK7ym7PEH7jtBpBuhGcApgZK36b10Rm9oZUu2JparVsQZvcANise4
/5UOB5jEFH2jyuEkqZF9f0DKIukuMSrC9+0jkpaxgBefmKb7OnKZvAHB61SIUsOa3UIKDLdTxF4b
5E1Odhod6bf74sopycblfiJoepGwE6ydlPX1xNYSKrpZv9U9v5pWPBX3MsC0VXqoQsM5PRifApzo
KGAOV8pQLhM/Q1yEKXMTOBliHG6qL0ry2HWh9lesR4pTKL2LT9n86lIX+YgzhOfYaLJ/mF/VW8Qm
U15QZD+OBYJMW6oHAuKzBIWJq0rg5sOYEP+DebNY4bXLjThyj2I8H/TiJPrxdkZ7JcBWVP5wOTrv
XbXYuSoA6bQAEP4rkJ50gdHi5vNeY0kcGWr+cdFwxpo53IxtzZBM8KAFi9RJFGVLETRcX7BjCzCb
bCZm8gzmc924jmXF73Km0H2fY7Bw1lNJyoGM+OGaCHCb81CV/WR1f0+4xIbeo+FjEZjXW216U3V5
spVvv0YYPCqo8T5d2OWmBwWjssjIQnvUNfqmolUyyJu2ZPD6bFUasR96ZVPiSjDSUW0a0Jhf7wDj
f39KhLATHLafNRtmLJouFm/7PwsCdIaHJ9hvxVrtg2rGPTeoIQ22kg9pJEETV8xS6ijFHL3DER9D
ebjO5uTJRIHW+omPeTicJpnZf9ZoI/It1jkhtyHCZ02EU2XhGrkRQdzv0kNPDUGurHrmwpCbKN7q
K5Bn6v7WuzuUiLobTNvgKFnUPnksmV0v4WaHsocQNyeqQtpzsXVjMMsyu+nB5x8ocZ7uoCQ9z3a8
C3cTAe3lt9dxR1nDSKd+QLApX3REIQV89BRSwBw44F/wrkGdiheRU9QdYsHjuIvnXg9M96pbq20R
Y4Hfm/II/YiNmshZpZ6fxHvyi/vpM2TRysYmGrBXPtgBSP7ftXe8qiuMsg/UkX3URnirMtJN2Phe
v0A2SYmFNt9GqltGB6vfa1SJ2lLTgCOeXSlAqmYLaiuQPR3i7kRkMjm/fC1CMMz1eN3rcipkkMy6
n7AtEbpLfn0J2Yj+1SbuzI7iPiBXjva1aSuLHuFzMwxRs52FQ9JdyoxhlfzjRNxmKhhfYDY0NXdq
zdTchPTxLS9vPCeoWoQPMuUYPSMq2A+BEhoI9kkJ7mS4ze46DqHU9dRRNFNVmObjDmbmuJ5PYYq6
AR7+n1nvYbgd98o2bnV8mYRQKOXQ08gzUuinSGnN0r2p042Zx9M4SwzTdFjK+94QGe4DCqSsNoSI
bY2IDKWem4VowTCuzAvkz/QpUhSJnd/P42G20LtaaZAa0kG/Nq6QfZ6VYf1/PWVZsXI9taPuq+gs
pvTaLKE2LzAL3c045qqE9mBk70u+0kI3MCyfmzwcrEwRUJ1THUsso5JP1k9UYI1PtG7ufepygRpS
HpW6d6ejsyYttwgEiME+BPzBHlKjKvuwk4CdAFplh/SrNDxQu5iKoTC+LP40+P4f+FPcExjGRYuB
1COhu2UFXzmLb6vKAWFIHa74VYT5OsG2WhoWUaKOFZaec9dsiN6NV2WOg0wUr6pBXH24mqf8Rzld
Q7/dfMmSlyfZHbQ+8nrT1V5tbqhdU1OxjDv47+0mEC4NDbMCglivfbdvmMtijQrr63FX56gLclPR
ag09iR1c3KB2EbSiP527bZ4gXVH0uVThbVVN+RWYMeBxaVcP5iGptdu/7mbnFA0pQhOLmedCKzLU
ung8QJbHxVsNeTIC7qfd7QJftvVUJvClLcqvrx86D/iJebwZLPw/0UTWGTCx/+LH8tt8aMPfL28d
GZ0cMBwijwdn7k8zFwY4JnC6U35Txz9nzQZwSQQG8+6xZPhYSOHlCB8QrqZo3uliMAYBKFV2y07f
lcop2Wmvvrp75RG4Gu1IkF/DaH7WlN6SeJJnlsjvsvx8c7qsFQNstVC+zFo2rI+vHLJMEL4lAlIJ
wUIBXPsQuL7BBgAaKV2N4qrjuzP1PdHXx2z5zh6qmdIdZwEh+ozft3D19BPfuoUJbCwL+1An46QZ
ctPFe/roz8h1aXu/wAcrFTpq4TahgKlx7J5tuLK//kcFW9hkEebDbiFFXDQCYtr0cIHg0OvLwFHA
AgLZlsX5Q5Km111T0tW+6qPhYpr/V0gVI7arFVKZ7SA81HWHFIPyFDoJG7H2ee8squ28JKEq5BgR
jU8/YxVdUGqSX296CtmJHSCikPunPQDSYTrsU++RLZSNKaq+vdyWVU6OwEwdyDeW1rz4gXT5vR/p
RH98nYXD4ZbHCU6u9EbuyyH3Q7dMG9Av5NeNuWKXe87T5g4zSzcATlLI6SGoB5dPsrTxunUPFakP
FWQOMJDAYYx7hw+VvaA6tMrWnBYHqVB5Hzh7pNflEEH+uQrjR5LOOHWP86zQCps2X/kkcfmPCgsT
3oP7OWcHYfeffwC2H8OFht0zp7ypSqWeJ1cc4b9WxB4FvQHsgpi0/ctRB44t0xbxuRLWj23GmZNY
xE0UXiLdtzKgQi2ALusuaDvT1wDgPjoJ/RvWA1WPlpPEwnJplcVe4iiKlHgnTkl3Po2M4T+TUtIR
d9LSXxFFz2SgbSQw+5FwmZXd7VqectJz0ImKG+9LfKD6+hKlw0rhkAiKzRLfXqTadfRkuVu7KmUQ
uGK+MP9h5dDWZfWTeW44q/npVglak34GT9loSvNqyqphALIculMDB0GLx2FZlviI2NGB/cwjETZM
dvZOCrGNg+Iq+L5sQYzBuvXBBMjQZcBS/+g7CZGe0UsAVjLqKhFUaaazeLj9vgTKsYmIutvXssVn
bFBkSKkwMsAGY5bdcITpHwbNSnmjvDrOrGviqniRmcKw/ea61HYEJUDlpGHp4jOmHjAKHhOD/hXz
ul++uaApHh1G9aswDcFK0aHcbh7bBQi2zmbfbNjZr3wCNIWqVVh1kOvGuqJNkwU15AIZdBExHKTA
9ihdghaecv16qZnnlcnG1TWT/wVms3etAL9YSFZr0HB0hEacxRmSp8rByDxT6da3HGCbaV2JAYKO
G3ZUmdYPWR7LayJSUn5jbCEvhTugW85fcO2BsmQtDtiC9OxsOXgtzFZ0wFbgPwYhYDqvFvqKRHlu
jMgSfrmlpBk/n7zGTA6fgtKH0iiAv8HVdYV8BzSfasEasELadRw5X/qosuIEsmiPjFHKkLR6EDyn
fstKnXv/HGFlSJJn5k707wefA7X+imG2AUlGLENvMiHTAkY2MoD5eW8Ot6zOxwyLMPY4Wc85zJim
+9Px50lp1123m8WFWS0B+W6u9oS8sWyNGNiB/hG6EhulgXadMLxORM0BaeAJvQT3ZNHF73KbdfWQ
gG/WbsNnZfk1pAJcLglFCn04LYGtmbmBwLo42ahcHlddcJ580UxPk726SljrevNrgB27WOJyzBHx
Nax42H7/HrL4caQLBwQn+b6u8jSNXSvx51ffSZ+LwzzUXBZkkyCFqitM12tRN5gAdFc+4KfjD9gK
Hdq6aFPHF4D99xrAIci559eAwUaNXIFl03jP021ssYEDRFt6L8CUjzBGsZd+bxQPO8AzdCel3wPd
/AdmkyupgQzbHhL35UEFOqvT5/TSkv/T8nxbnLRtf88uS33qMvPUvOzTGUqHSXLDAiIuqY7A8Z+d
itJi6oP8oT5ncMFTyD2ejP91bJYrQTK0kGN6+8huZD4+nNcq0siB+G9ii/N3wcXnCZA6LdW6k7IL
SgfpHCxICNpoOcK2kQCWCw5KsQAhjxDGkCiJjlcCvThIQVYm5yENVsoqQhzjQy0R2s27B0zHQiaL
uKKsKz4AjCLmtQkPsxzJIrrFuVGOn2p75G9qmq/O29JIw9OgGje78NJC6uFgI8jGLWIzQ30a278p
vxj/nVN8c+yBAKMpUMKtbpgGc/VQyhE0FhXf4yUFiVAJY8BGzypCl7Xd5bgu9Nr3ORg32Wp3GIc+
8SBt3hW1uuwrnqGiUTYCvA53krCAkDWw0hXvQp8K8l1KAw/CGf32CPEwKa3n6oFU80M24lVZsm+G
aGfoTAXq5+oMwW6PjiM+eDUkOQ4ooI0sJ17/xtqoIZt/vGBNpi6HfF3ApDbzNYCkv/fdW20+dTu/
PrWjNYhZL3rrapxZj1V4QlJwKeKQbA9q25DGMBAzyOQoQ++nGOm+Q1lfc5KEW5B5NAwyv7SAZ0vY
B9c7nYI9gvSn2CRqmARWvKmNR3BEFO5B1ynQ+NGOuNZWufmLi86W4jO23NAtz7/sgTMgVoSd4uZV
XnnIbSv0n63k9VHY3qiZ35hUzxQe3rjyd1rMyLvoBevTfvsI3kVbW150U5dHVU9iaRQkvMcYnD4k
dlym+Ihgh45ruSXjHATBqfF+igEnutZ87QmuNKknzSU65wLsgGVYACGoVt20b1SYFOXRXEz0bJ9Q
u6i/JGIG+6F4uNHG4kpXPHKQP85d6M32P9Q6xgCCzUwKSRPi9zkPlN1AVwB5PCBTe3AhMDmCa0wS
5syNcMBOCL1feCcIBR/co/a22yoHSSmrbKV6mHbgyUO/BDVLFX9qxUZf/AXF8+xvbBh99fxs18vh
uhHR04HhT/o7Ma4eLbDWoZx6LSEgdy8ngWNXcOGZlBx71B2iW6sugUjvlF3mG/M1AHG+xnn92P27
jFPCa+zw60CFDmbdpF3aS2Iw72BKWtjoJdw3ndndJSECPkUp8OBQI3t6MLO/Uw0djUzoYi4R3Jzo
OyME4bzjLLH2RlWrjBy/tcCgXun4n5FbgfU92Pyh95p36siO8d1q9cqFDZCYFwCKpaeYeHmhEXGS
dN+INTPduCQ51C1oEEeIDacg6S8m0R8352GjQ0r7UtvSAe+WZbciT0KaMdo+GgnWHIbyOIlqkDMB
p3JDmnfJ/YAQso3wE+WCl7QatYvFJFrZjdJXlYWwADFzsGRDcSJKYu+dWBCLhHAYLUF9oIRZT/Z4
mHJ4hdu1rZKWA01j9sONMv8mwBsBwgFIiUebhr7+vYuhGKLCd8ZnN3qUbV6bmoJcviKZqN0hPXfN
FZnWQaEom6oIXsMA6PGhND9bSwJrOKZs5WEFHP+Ka0WU8TsPu4B+XYdSeRfIhPE1x78X5UFqLAOv
CtW5Fy+f05h3TBSutO0LpV8NJNf1XOPzndhmS88jVIzObvKO03XfsFIw7ewGscvTsx22GepSdkc9
zp0a0cPGZ5lNhgVup1csNU1btq8JtAHa8AK86qjRTg/jlE5bDdwJhFKKEpnT8IPMzWoP9gkqjjfE
ZZgNXoTXTtuZqpSOVqiJd1IYmNXI3f2yGfg2nxo+MK6AXF/4grVjoHsGbVkg6Q0I5dfPKl9KNF5K
5KKqmWVouEtVtnIJ8YVZaUD24szdTSx48RCKL3r8xiNMQjQlabPfucMBY8ofHuX2HqWTCh2CFFde
dVKIwI6kHVekjGxE34BkS7iJtb3neBwsvy2d8T9EUETjdgL7ndZGM2RqV4KewvZreY+JxzCipX5x
ufP3XfFdZJ1l/cAWOy6oGhdnTYLX3CbZqPz+vQ3DiBexvRGGjxAkFNh8Npn4UzQI6hPCvz3d3zqm
w3OYxSWn223HCh7R4ivtHasnu+0OEJj1inkDrsHzcqtNYB9cg2+c9Yo4bP3as8gYk4q6cwwGjbCd
GCFW3Ixe43vXSPDQz4K/d0PKpiPluILCWEM0GdWTG6ECDu8O2ThJTnEozAQJgTHMA1admULMA19l
D+YnH5yEhTjsTELox0qTzuyp3KQ8NqVrS/bhO2k5BsTkgkJCLy1r+WXLlJ9oVUHI3lTbUHj6zmli
20m/QFV8DV1xGGiTGketKfU54joKk/ppWug828lvdU7/m7JdLHKjn+4rIAKyIOGYwCYda92tg+fr
fPp/dZk2NV6QnwASdAYn4fny46rx20UlCorzngrQLh0CsH9HE5EjYVMtKBnqSxTV8j+ymCjaLXMx
56YRBZTuV+hbgHetYtdyBP8wLFEl+TX0+cQf70b/3Qp0sS21qVV+aJVzlahuD7L4t+jM0dMZD+50
RPIi5vYAB7g+jVe5D+1LBboqvlTV3mNiR4VC4qAxZKUU7mIe6bamVGWqGgKyuGtU8IWby6MJikne
52bZokbaph56eMI94i5iXocqO5zStIB0Yd81LxsImglpkwzWV3966nm0MBGzNfM9RPcJ9n7HoMQS
I81OuYZ9NHjngJGovuSF3fTvoDuK8lutzFDBMqGBT2GKjPxFj/vY4hpSOIRNquMXBWXtZa8qkDR7
90U+to3v8SeXyfqFE/qdBjyr3g0FPinbExFA9OPggSSSn/RfgZiqx28x1TLN6l+mxldxic2lKTIq
0YDIYuGo5zinyo2WrYT1YtMv/6gBrOty5Rc8rImKLFnHm2/aKB0ozSIOWiJce+MMQQmydpF/oUmR
5dOq77lT8+dNjItNdJTlY7TmVH33g7DJxRYMqiSWdHcRcNLRFrEUk1VGxm8OqRf056YDGcjWa6az
BjBiKQtcIpehD+bALo3JaU0ypuDdp/3huk3LCIclEL1CTJkv0wZjn9S0rMRHznfdoWrnjlgdDw9i
OxOcTt9V4a6DFuxaD6oXafQ6JtocBQPzr3wvEJMlrl0+KXKm0pFiN/Q8gvVSAoW4jSconQs2+j0Z
bFw7u2gX5SiJ/MlXfe4ZTHHLnygRpN0b0MFCbun/dUmi0MXWmo7mXnTBrZ7/ZVuC5Jbr5YOd27+p
xlZ6s5eMMaVdGmsOCAi5n4SJwofIo7X1Y8kjgoDCZ0Bq+sMcFi+eal+bT2RXDIp5lgkK+5OfFaGv
oYhqmLaRaQ25+XC2ubzydAiJK44I7x/+glzVIZItq3m9q9ZfOQZZuQ1ns+/gvy+OOT/bLKNadstB
FuybMSLU9mxiHfxTnwysXpCxVcg8gEXPP8Axv4ke1SBID/EOJfcj6Mo3DvgX1ObMgicGoBMtDt/Y
/PXnr2K2sLbtDFw592RL9VYTTEbmXB3vSECA1CCmyTFL3AAHwf5PwkdkntxRKlmNTsh0uVVoFuW7
tYy1cvRBoiMs5AK3A7yWGfyVolumV/TM9/Tj4maMZlT9sIyc6C9TqBg944+/90Zy/9N30jgBn9BN
J6VR7OtmCwsTui5lT9/Mq/Lpe5npNX9fqd55c7iQAd6ppRHp1Nq+Cyl1iKgl5QNNt+Ov8zGtvXGB
tSFoWGfBFA5J7OLqjTnORz/JOBos16RFw4blTC3cevF/WtAdcUysx/7kB+B/XVjM89l20FnQu0SD
pdOE1kA0SAxlTwBZkRDYCW8EHdirsXGl9P1JsyRICIo49ghAVZvA6TfEfX42YDDxqyf3lqF/j12M
nXwR+2RaCrbGD9SJ3oYJ3fXegLiaDp6YFjddveotg8BdeCgK6KG18BsauPaC6HY6hTEiySO8EEtq
GV687fXMBqeTM2Kv2LV1uB/cCmY+ffiVMTYVGJ9lqhk2kgiDYZWsQGmcvG41dMNEb6T/5basolyc
qnX08I49vBsGlMsHUS5unwtqk3yNooY2qe1fi/Nw/okHaOPsfNC7WIfibxSmsnKwa4Yc4+WH9ouJ
Iy/ONesjHMVo32i8InAUTxmIhzZ2xk02IA78BjTbK4sv76ZHInKo35Mlxo/sdURZ7NnSLRWS5Meh
gvA1esV3chKEl/GwjXI/zThaxPJ9zDG7jtt5hjKabQ4rTmGJTOLpt6Ylx3ELKH94/s+tSntCHhgp
+NaRA1EdnavjuDuEh1PBUwjqgk+oPoU0v1ZEGdNuRfH4xfB0b6m9GMeChEUL+UxF7pkGuApmYVQj
glAfJwyEpNyPuwzHbl9NuJIansYXR8Gp0gIiYjn3isp8RjrP7HT0dRPE2pWfa0rCWqUWzKoGNehE
Aa2RhzAXya8Nver5l2Dzm7m76XLQdcrRGD7xoCdEwgTmOnjWDp+otcbJAJFA1ALhlNRIMS0ylUcY
5+LVkZHv/MLK1lMdjGvgibulrWcovzVnN6L1fockiIUxWHnnVKwc3ZARnmLRa4tJaqB3k3Du7GL6
U/RtUKThxRTDAPiw9BuzAKl6VQADePN49HvY6cmxpeGxoZt7ZSvIadkkyRjfvWVzWQ9kBb3Kg3HV
0HlqqVamhLI5t2iSzTZHahbIf2eZN02vbBrK9+ccUCLznV+WsBCZJDwZnDVWxVWY5QhSn/tIDhxX
+mm2EvDWXLBzU5EJKlJrBTGU0xbkCqmZ3t4MU0CsCdnF6qjXrDTTaeJUyT+xcatqNdhrhCBaLn5x
LiztUyhK+Z0aMJwAHVIFUU23KAiQpqqpNydfwxFgSkUWxLW5mYIdBSkdcsokMMvpbYtJfd+b0NW+
+eh+D8y9HRUXAOeRmVds6cQaY13KdUzYIcOOuUmcqM+eMPrzTyFM2rP0dRMx3ZXDGuKKK1tryvzU
NmE3y2+w/ppwIu6u2MsnJLvdy39BnQCBWFLbjp7CYWmAIOcWQeekvibeJbw7Swb/dvPn2/Dj2LgQ
Ca7tVaKWfA21Uj2HAopwIpYaCq7SOTjfmSIGGBzDXTFXjY+f/Ps909sob1xW08Nsqb3UgPGrvtAc
nZdvhHuQPbu9h9hhwCj5rEjHRIk76vtqjX+iffFl6t/cGqQ4I+Fmt9mX/LJviUU3ohylAFIL0PYy
gWRCz8HiQAsCqkJwwrKVXvxV/mXdfwEpKiIsJyrBCdC70vzjanId+sKyTARe+cscNFtMbJXXqf1W
WOuhkW4taF/mBhqvFbgp26MOu/BDjs8+UplJd/k5oYgP5dxg5Gy9beHiI8c3QD608xgs/eeIbCB8
Jzb1J1JsECFHabh7q9qtdDKQieG5BidghPEJbP+umokEkjupG5dpnacYSo4bc59usWfVUoZhkjBo
hlkNHKxw5FI6jufhzO8hw+OTKZEl9fIWakDjmsQRzTDR3Ox8PSZ4mBSPtOA9MVolOY2SAz05mCjY
rRvBS+mxYFGC7hdH5Hqwe/Kg51sI194We0voUjILBnqWgN/ssQKxz4zXSZF7Ez3l891qSDNLBOCP
BO0wxrxTiVPkZn4AM34W3uB1FV97kH8g08k4wBiENAEsd2LV6E6/ZJxugKxKcdmXXVU/XK+3ZeoI
INX5GFMN6D8R2vsv/OsxHauom5b9aWIcd5LjNMkachFM7SnzyvlFldak0cfEFOfLERzIgyivis7c
Pbm/35CRt7uD7jTExqfJisNCaTllnzhmvyvB78Fr87XpEZgJli76wxILNfQcF6Q+d9dhcy1yFu06
vx9lE9gU5tO2HFQDcIpOLKSw4Rul0sNxRlHRe2BuTaZl/ucPF1FdKaknibdRf8dbrGD29GpSjXR7
t98GKfIlLD5MP39iGZEl71nkOS1KbULaG9mh/HQHUdUtmkYHsRxbInJH0Bvpzh+PPFmhGrtIzGo6
67aqxyIanmus58UVzyDPgre6zkOdg27bQapP8PtbUzjMtA9RDskhAXe1SZ8AaQH8uOO+U7iasOh8
gQy03cp/dhKfprlSv3KMyQCSLgNvHnvQ7UgN1IZiaw6vXADhFJYuV1rR6lw9yd9mkRwv5w7RsyY3
wkO7dUzxlqFlscxg8VdpRKbFcAVX1J36bN5MQC7qVTUOAE8fJ/7XIK0LQWrSxEJwwDBrm9JDCeRT
mDsc2r8SiUZnqZSwOHccw4UToWEQa+YoQ6XUPEXNAd0ox5c1TaaoXyw4Wo7N3tesGQDzW7jlkzYx
2X9UIukreWI6/hMgy8Na4/dFn7DKgonkqwHUgaWLZhaAR+qEVJHW2wmzvNysgtn+/XhOIeaBFz6T
Iyq2Fpb2EJugyywUssP2uwIcabiK8gTmpGOyLqEUVy1ybBPWFkSctoidxNLD2wcltGexE3060D5p
SoNpPqAjaWcqCYeuPnnfe6R/1JOhdRZ8OjgioioWx1FY8dNs/FgExnq9YoA33bo203366/gV0KWE
Q5mK8+mQQNU7B4MSh5LlYC4ZU6+ng6aP1qCujVnPH61yorqMMYrGVz2kgmSDycFsRi2GrijyQers
YXxmFKIwW4HXhjvXxm5YqKRloawlMK9dRCORfY//DG55xvIeThfnFG5l1/G2sRG4V2wH0KE+Bp3R
3eaX5Hub7mCPn1EUZsK3GUC1RS1vRj1EpROg+RZhj9nbXNc7Yig7FyAT5WEZtTcAx1mIsPC/AuIc
rqzi1orpcVh8ZkoMYxl3q/9N63IUPTcZC9JGPJ24MINPT7Lmo+gmNHmHzUrbR1gKKPbkNeUWlCMY
baPSfe0dkIPJH6+B6aIn9sb3+/N/wHN0FgvmRJ7bERepB4x0YAbGI7OYDl3dYhuHbZq1IUDKRIoQ
7tqe+dl/UFA/aLZuKW9ZQ7iZfIEd/DjXyS98Lsps9rzbFkYnW6istrqCop1fX8sA3bN4uMWdyXeE
0hVg4S8SGlWnRDXmiOoTNZDweSaFf9xFwr9WVrrdsHMbCSRjkNN2b7ZXTQWFjZZ4IzDB8CapANXF
iaVnMttl4FCvsY8YJPdBO+lUC0sl4GkmKS12YizkEo/7tfDwY+6O7m5P1QXAkd/QfrKMgT8XMSXN
cMmoRmom17+4gjgLspL5pr/xluPR0y335/kUu1xWGbAtwVz9zV47KcWOk+nujOoiV46bnckJmWc4
ZzINLjmJ+cH2KffPRs8jnVx34EYzTsMF/6i5fWZTx0jpE1errRqw+tccKXiIc3YicaBAlYLjri1Z
HTOkmUrrc8AEfdJHpDxriB6/uKGLJsHZrgK9uZ2sQSEjWRPH4HYlZLtUucwHm/dIecKlCbyf6nOU
zqH1l+mBydAbq7kyZApk1Ix94RF4C3PyypGmUxr97PhI9moikHG6/HAzamXNvasMxmpZcnnbkQzG
jKieQWaaTebvP0raF4SLbytrjX/gTqRaWN4FSXVTcrMEPyH+mNaiQQgfTEtvcbHuP5O2D895z/OD
pzSOIWptiiv/MguMdHF5dwm2ks3O7WKYKaCeXXWXwy6lSYc3VB26Xuq+t3AC/avQTTSmBaOSwz7T
Ib1zpvjc+V201p2Hae/QoDCYXHoITKYbU3GRofkHz1oCWqcWXjMFNcAB0qZG6Th7+O8HZQgiTm2u
F53ONJSYuITeQNYL4klXcNcGUF9FLzCaTb5vr1yl/8SVk/DuvFL0P+lpycA3GMVeBl8GdfxeruHu
yYzKNGL9Sq21X8+/vxmm5mvoHI7FlYg/e5tp6dileJdHzQlacVeKff8yKmWD74YxcYVOzesYRiYS
EbR3PydGiSa1DXEtsHeqo7Snd8KzIyU/ZFS/hRVHCcYR62cgbtfvGr3OU2b9eW+KVMO9JKlepVF6
N/tjbipP7RxynR3ZOTfyExVydb2SA3ikRaBCna+1e5crmn6AafBlhgS93Y+BM93D4n8IYoIYTks6
B5794f9wddGMxUWW29Y6KRGROWonRTSfYqEQZrqG8MrvRBtw+FmRPPOYS9Gwc4BDzw7MJPoHKCPL
Vf7UewPUMkUXYBRYD054gTjhAT1fQq/BzW15Aiu6L1dgErqRQoSRBD/YS+QICWQC/1HW61Sm80vc
Zt2GFlvq8lQSWEH/1BEo5+0bXZoZeEyoJWt1EIzWqVK5zvvUmetmmnb4/2Zs1NY/WpmQeDA7BCCc
YnvjQdYsADyDD+SlLRBPteF1AZavRsCxYK/WMM+1/eoP3ZLbbgE7mL64VPRD5KTK7MfuPDK0QSSo
bfVKRdmqeHR+1QjOWinG1XQOUrIyJH8+4xNMhH6AIDgCu6/ktrkTVmLhsN0/oTg73dK1YDQXft70
tuDwq+zSFzIOxiRWCy/A6hVff6XRri/dpZJFftKkQ8Uyr8XbhT69ibO//ObUu6aoq3/Vuh0EK5HM
oiVYsoQ+ylEiKSjQ06u30n+KEH/wTFnAsVlJ41DQWP1G+2QuUhJXj3gLwpINpOZUBptM02cxywaf
A9/WaWoU4Pva/aTwRUdvfinO7Z8eU4fitkAhqggTQXQr3kS08/Z9sw1Tzjn2kQFzQasY9B6/G/7H
IL/KXJuGimwRKT/GArJjo5NcCtJvINBuEwW6WBZaKuZ57gLQlPdvRCAHqqoVSgbJVNYVj64aEihR
2tAO4x2vBoQPjynZXu2CftMmHC4VJMsxvaZFhNJLQRCNECzCsUcFhkEY13tq/lnYDwXzeefUpR5l
g/GD9YHNxrxNXyCVDT2Mp4/sgxaPw2/zdunI0eSaZ9Tue4BkHPRZy9Ctj0+qLYfLN+NCY9s1T9hD
uTN57X2s1OHJVUakWwLrvLW9fqxRE75IZt9ykokU9mZrqIfCdcv21kr6DQ4jLHgYXDoaBRuBYKC6
xX43CrtQvf6gP6i6hUrIIRWBccwSe2EkkhGc1iefjrRhw0p/pbVa1zgu13tkDfC9+daqzk6QJnQS
ShLAg43Ei2gDAqcbVnO06GK+FKsckyvXv7SPiMGsQpwhu+CPVVwBt8Vkqdccjko384299dsxb+yt
HCaUE00+BTR9fCVH+8nBa26OkUnhaMLyuH67FzuAN346S/Nf9NiX8SQlcixoGzTdwJzbByMfBVLb
R6HGlhAln3EQe1D52L4X+6O9zIBJtM71v3mjHgN/NhdieCYejcG8Morr6Z82CpipzJQTUHn0ciwl
1NvpzZvI5AAgzKQCmwWoKOUBNlmcFHivGhyNiG7f6DCUbbuWVz/HJRZVEz7yGLSd6n4h7I6cSwg5
J4f3bwB3ECj+8BxWoQsql0Y3nhQqKU/a+d2jxFAOYXfVGSlE8lFgn/H9H2PU1i45E6gin1qMVu2U
NwdBGD7qqvgc3PL+T7sOwQagWtg5axuiwYWWbEQP9nmZEttATJes+ai26g3oK/MJViHdQylKv+4X
DglbRfYK8NVx6jsp/D9ZbU9jc5H4TY9ujuN8L4OtoieiZWa0fp7gu4F8DEL8qJP74aJ8vu2XTtHU
xofROi7qTSdDaYlmPCWmcFUrdJ6JbcLXq+Xkfq83rcTHdXgcpssLP/VGAWCkEJnP2RIexxJ5DqXx
/XCXOrwVfl6dqnEt/rFQxTW9OwSVKT2NX6m2Zl0773RuA/rc4D9b2ZRg6jSTPxePZMnWXUp+HJYu
TNiW/Kd3KB8duyYI1tP69GMRFbZVjMzN2SgxaDwpo8hHKAUWtLXsvL5QbSnKyxso+hzMSDWwpMZl
CU9JYMve5HK0Bwa7Xn9v8QqX7TQbEiykiFCwIC7nDSfqmUyHYFDdCk2ZEYRMEzZQmFnQksLQDfZy
Bn7N3Lv2g8RolYfTRLMJyiVVKaGev8vULd4H4rggIjgDDUbOIvoQHHU7JfB27hLDJSzzZfmGVd9x
NXLDaKq1BWH4ZvhdUhZV0d/LsFdyiqRK+4/JWmMo9VhldqDEuPMvl+1MW6R7GrLoiniabxO2Wau+
5qTgjYHCMSBu/yveCkMB9pUHsDwfkppFTA4OKFrLRDoHcXGGRZjCuhdSN66Il5SQOFL0yscAHUyD
zoTPyx//Tu9yeuhG2bIQPDFd9zzGuY6UE+JymNJSmr2/fUkPjW67hWzpqjRrJN7dJpZwlcknYjt3
da0wZo+3pl5DxcSqJOGCFJoKwK5dZ2MZ09rswjO+KtTGTWzDFVOVr5QtlV5fIAsPkE8H+E7exe/T
KhziW++Czxolt+Cc95M4szrMdZVG+S5ZPX4dES0nASAoymbwPsKUQxWeuNRLzjG/yP5bKMuFE20V
OnFKJTgO2/Vrk045SW4ZA2yIHG63fbLsqzLqPnw2zF1hdqi8K/niLEUy70nh+Bx45TKO0gOTCe6W
swaS6xZgIlR3miAurdEnqt56KpqrUgmdIVRKd14/BlCkO3wbgTqiUch62sEx8wkIxawmO7UR2atZ
l+fIlqm3A1j/jRMxQCngNKyWbkDmJLgTPDFszcdAdWdOre0qoCnH/YkyiocaztttQUJdBzd0MMA1
3ktTprRL0sNWbgMdUVz4tSs7Zy8nMpiy6fOtBDWN1vIQhcupfmpJ3OytMQCsJ3qQuzsJiqFZTykF
FUv1WJCsm/+BBUoTu8hXZudets8mVCERXhT6Tn0/ty4qfYjqJbT95C/4KH3SgxzLoH9kI4x7iouM
SFSOvk1nTiPXPSghDpkAc+IkNN+dWcDP7Mqj2HAJ9U648WgakNFOIdbvUSHod/hDCKyM6UZWMMDb
v7nfddEo0FTdPofWfZGY0Ngt2f+g1cpdVUPokSDO04xjsgoxhtuTEQHGlIIYSL2JzJHzkI3/wvQ4
pa7LxFi1LT5Fm7FLJOV2duGa/Nj+I44N7lnUexMhbgmV0qxCYISH3Y7M/lQidXk5ZiuzJtBPvzSZ
RGgvaySUsRfnciorS1F76Vu7XradpSYTwcwN4EH87+wZ3GNMRULdrtCsoUsaYW1b3Moc0TqkRdZ9
MIUl7AD1HDJse+iXBzx1jhbAW4GEWn0XJ/+lMdxL2ZCkOEKIxA92FCloGAC2xxyICqa8LMNRNuhG
F0tYCwKe8/m2UZPL/D69gRzOh7ThfaAFHUOX7altZZ4KgKCKAWCFGJphWfTWM3aur5ajlk8/YwKu
jEjrU21KIvWt8uab/qyB1lJzifNLgDTAuuec4sLkxJe9OIIKcZVqLVf69H1VK5poYVFsayIgPs72
ERXDNin7nROXAGpjHUzIYajjdB9uKXyVH9E5pZ5EPxJZ+QUC/SdICj86PMshhoMsK4yvNWu3c9gG
Pi59al+50k+lO9uCTUIlVvlILx7fVhvGYKhD1ubouN5ngJN/L/rLUHRpUQiRVmEcZw+Er6mxAs6G
VMfCKvwO/J943foF8P5J9Oc6Y7WMsqJzvfF/55GMfe5gwoKDz+WMk2ApwJz7TIaGedB8JeY5uZz7
CDDRbbkYuuzj+83h+mOneJGUcK7KWiR2wxqTbp4L48Cfdje5cWVnjerMlhx9UMeWEbEKJxZ6vj9V
10jI+WdLE0L2jI4h3HLPzeSdzRcW78jfOsxyExkqPsY/4k5xs77k9jrfa1rtidGegYzW9C2q8XOe
P36mfUR77GHbJdt9F5x4R25Y162sFHeoMebjCvO3eJUtXYWEiCGqtuHkGqDKKDgbt7bUA4tI0RkX
0jjyIFyzTfi43KA01+0XZPOc40xTYxkI+15owDDbkyXqfM3POAxlXs2HN8gn9C9XCRAkWgtOpLXA
dGoMkpQNnmOpgNMQnarfOqo+D35KVpxYL4JWe2XtPKCbL12ApEIHqusxaDkz8iKwJPdj/ieqEepE
UsuPVgN/H8nrkQKzglXUgO/LmmPitW3RJGngNU96dyqUzxv3fGxvJsI0dq59r37u9PczFiPlVDSY
D1mUjfmU/r83jtXbddma51HfQ4ty9mgrYxV89QKMJ8beVjY07BDMVKrOsykC3V+GU/qENiWaaGzO
tr/Cm0tAjkJRJ8hKTY6YQVI+/dP1urQCipyzizMFYkNwKL6RyujVfeUU2FnLlfBSyGwqfyIpaAJI
z93mlt+RiBCadzukfmsM54G81yp635qBTIC8AlS4bymKpn2iLoMriYlbaCSZVcDvuUi7JzW6Pwga
/hvcWJ+sZPMUnbyxqA+kiPUN7yC4RsizbbIBf2vavMusXqvwMf9iIOvYbwBeTLE2U+3RbucXBxHS
4cLPBiucVNOQDmdkv3GRlxn1t5ROAjXVG9/uYK9GCfLjfKAxk7fEvG7KySQB6+r65sapvXRMbRsD
8RGXXoD8UAIFBQ8GoMZajPR84GEoG3r1HvKo1c7viF+yfJx9bL0jYL6Qa6lBH/YqVjfbpq8IDyJ7
0i0zJ6dsTQjdWdSvw9afLzop7YRTVaSEwl0CY68JXZ6RPFJ0Zxuzzy9m/IdV8Npb6jia3fx/3qpu
/VUhZdlQvLd5fIR8f69ufxvcRemNq+f07MGyrkrQfpEHQ2crJeMciRpGOJEpVVpDIi2zezG92rJN
Y/g9KbXNhytiiNmAhH3BjMyYLX6e4ncebggifQeGb4Nhc1RX2MGACDVAww+YZORnIsG4jA6nYo0E
TCLEwfEbkLPUBK0RnRaUVIpPVwklGD9WyAAnbwNpJb/SGGvPeKWiY19zJ7Nh2YjTCgrFl1SgShbD
DQ8qKLbHp3BAkXN8GGXmXReeEM4yLVj4xvzdRAI4+wScNUBcvT4xaL7mMjlIbCOhUtvUElMd0604
kWIejuZCbPIeN7iwApfIqHSFe+HvxJLnn7tnZL00kEI88lxxv/AGOsQVLKsy2GEViMrL5T/jCPwY
e3kCKtvCM0LcuMEVFhmeM0SYW/oO5N3KQK+AafyDoe1ZwlEMc1b3+tv/GqyvujZJ1mEc3wPNUMYG
1Sky918Jvn547CEL4Barhb1ZxZvvCYWxUw+4Th//qzuEb2FJTCxPtWPDv3aBMzZzdX4ZKtVIH/Ps
JAzMyfhGULbVzN2/bJYozAokwvbmB05iu3133HBdksZJk625kGC0eumOcJKmhUFT90qrIQruewTt
q+JaIE7TW604xtaZ0Aa4KJFkLvV0zvKCxFVFqCH/8J9n586ygctqVDNOihMCmhqtzaE9GPTLSdzl
XRgCZ3MXOzFCK6/lW5w9sbPkuTGxKujRl1YuC8/Ida9+P5Gp6iaejykDN/FNmaK6CqvdAalofFeQ
s2xff0pooKX8aZ1Ezo6yrIWTyU/gSg8hpYWbupXQkSsgNGRACM5JLD6D4TQMyHnQ7cLxpqaGOQ+D
1HRyfUaQT+re3JvCo1CaSMoVZAbSQpt7YUZuiAEhEtzmGCf89NxMglW2wWqY722GyYnd+ZIO2/2D
lDJbA6pHlL+wN2fad0CyoEw3vRPY8hWjyvdu9Dp6d2n//94fsBR4gRLdf2dSYon6Io8rp4FEqAbo
mzVb+zNpTs4e79XGx50p9kOnuXhaimKRYSskyPfA4aAA3hztGYLMUyvsilWw4qtl8ltB+Yt6IZMW
ESzuQFQc75Pfn8NaTI/HxUUWVHYMIyDuJL2r0IsG4s6fZxz36F3br6sE93OTzzlhtV/izOUukq+V
oqZnwqfo9XzYRH94bi0GBUNEN/ThqfAj0kJGWWEEkGzSDaz50SgGW7i+wDyHB0JbuQhZ5nvWNWMd
dR8dHdAxtmdFWWttmWkgt2RRxhVAcZhkxCWQhXi0NVDqYJwCd/ntyyKkWjrWwdQx5qfGv49pPWS0
bAMG9vkiFZQqmc2gtJGEuheRUt9n6H8mLMW6Ca1fmc04ZseBGwF3dCrWdr1hNPoZNiMIpfas8lEp
sL3/7lmCFTDPY5l2Jyy8NowbesQIkbzqvajBhZfB5pECDBIJBqABycvz2FfnsNd9HD7LlCmWX+Nu
S5hGAeRkcudyZUeoYIVXsFYl9HmfCfkUiFBnpCtYXBgWzgVcf+zj1Vz605/GS3KGxCc8RHoP72CN
JJzrWECSQSykb6t4wH7aRkw+OiSSeyoH/mBL+lFFAFIaXql263bw9Zy/Pns3zrWoeqey+b6esXuo
h1UHQMbHuLLqf6NJvhR2S81DA2ePaRble8oDuriVLaLkF6b3M/yLlweDUaXqtGuD4R/2Cs8obUdm
4IqZe4UpQL0g0Lu6PA2ISwqUFthOIANqijVb81HvZAVh8Lz/aNM10pfdAjn/z8do4VSfIMAy0Dse
5/mKAElUPz0a64lbImiMqnuFYhFZ+jUrdkvvR8iME1Lvw6Zy4FG+JOmPXhO0Z6pXbFL6OWCSTe1H
XQFcLSf8XdAfoj4lxGSGG+e9HNYQUnwf33Rq8iuQZhdRUaVluqu8ORLu+y6c0vpgnyChl8DA53zr
HP3kqHWQHmEApzxS7YomStafH/eQD10+ncP9GGI+NOLKvo628yG24zi4iTgO9YzMoB53ueU28bS1
5t43VMid3yQsgTWYfD1JdLYqmaShI+iRmIu/Hxet9iLSlz++2FtrklQGGRKb+TTyztF4YTJrPKRB
4j4kvFH25w1Vm++pCvKZYV1NzMwOctvUaXbbwtiFog6m+1LlTcicGQG6MRN/05KwDjwn+Y1jyHH/
QZL29jFBeb57YVil4eBAX7T6jnlHBpSdBA4VwWZuxsjGulR5FnUXnHpyNKpnF1xciZZ3r5t4b4ls
XoMaB02RTO2jdPiRBt6FSbvbZw+Y4pdx9S0nZmJzkqpLySQaaljvLBtUo6ZIDkanOBGjRqtajjcg
YXxT1jpqORLM7mqqPb+ezmDkOx4rlRYLi25yd42gGPdxM/rDvCue35rRcDdWbfvD06CH1r1FK0NE
wBUaWUe1uITYfNNVLkVnu8oHYNRRKc7d0Htrya8GLqVd8ci3oA85wYJTTzq3bkVu3kD/xtt5hpiL
yhJBnY3Jme/J6AZNWYIJMa8AuUQ2Rq8AI3LBI+oMUKLHrn/WlOnsRDQj4efTTV5632G7SSnvzjtV
7CaukKhAMn2EvIE6T2GSWXtFeYe8SkmMUcwv0oGMpyJ9YFLWwu7kYL8gZ5FEDFLyAY9os6282VZj
NfJngTKTrgshKakV+lwg3bmmxXV6torAa5dnU+CG8km36OHNpe6Hfw1gpjmHKOyibvBaqAsPoYCD
Rsw836hFivK9EVrDJKhrFW7KbTp4OgBoI/TBGL3+aH01XDxQOBn1wQy4Y0aneUq3NXKyNoNE4K05
Wg4p0XawsZ5SSpLrWvprQ1/lZhoy1YnJEVYLKnie+QoX/qC5YQ16yhwDBvUCqKpLgnp0wDbAkVq9
WUU+26TDpJ11JQDVS3Qcxp0kiOkf5fs4YEW1AW1BFSjloC4hRFglyXEZoNbnu6Sihq4NazMZgCiG
ISF1JWtxcCFXdHXMZKRe+Mo1FADLyTZeOFb3SAxOYKDp6k4tb6XW+s0Q17T2rfbyfsty0wm5RKRP
fyYeWw4cEXsdNLWgYzOhH2v9Wt8GXz2GjKlQ0CRTYCfIs6sPHBdZe4tOioGSBviL8FsafGLLQy5U
ybt3LpOH964tQNWtA9JqO/OjEvdd3hb5l6cpXAk3oFkI+AO5S4ZRTPiIAplqesGMD2Ar4dilsm0P
yZ9/Gwx1NeXXOfjsmTbb8vxVaZzUVQudl79J9RkEzRv+WZINly3+EOF8YThaH4EvOFWxiI7+SyMc
osPoTX0KO7Sb+af4sev2qGd4IfPqMgiuTZFL+YU2CkJoO2H4U8RGn2/W3l7FJ24ztUOsQL6FVspc
aaqOCvWy3zoEwAiWUiakkxL2m79LG2b0nQDBw4lBFNi476gk8IYqVl4tC34wf3LsAzEUoGVbIfaD
8KawqM29+Zl+XZqukvpc2N743MDLcm92mPOCnXgibUviV4FdWMMIDcfKgU6KZb2xbD1CcK2otLGs
RdftVsMlWgoDUg4tae7f+v3g3UGToZsQImSmjDyoYwWBwNtalSBEsjPX6rEvaeNGc5jUylxv5a8C
pXA3gXTLhOc3gbQEPrQPDTn7OjrZYpE6/4e9I15BjZV2NEU1wPdTsWaNVnTtDV2/nHvTnDqphP49
wF6XNdVatGyYkvFiJtDq7CLxZWL9dYjonLSnfAZZZOjnt2iytRmhD2x00QGa0UfbT22u0j/8JWDH
pHeEt+fd/MCAjsJ8qyOTTjvNBC+I1dz5yWOzJn9+xfuAQCgYBXIs92/uHyxquoLx2mHOt0zQqTus
6tZPC4qpNQ88H9l0cDTGKMdHgQ0ZHyENbelILFkx9MohxaeG6sXV/xnVYhtFdHHJ0lHkenubYbjq
xdfMTw5HCkOglgYcAaWCf3wpvd3J+7yIVYrMYxrGFB5XquD2hp4C86SNYaf/TJK3w8QbWYZ43CNH
AR6rnvz5VVZSUO//cANoFCuRKiG4GyNunDhwF6q12LilYa9pDptUYv86lbq+zpSfDSjh8sfsCkXo
APkN+bYZ4Bh/Xqhf7zSiR8sHE995JfFnnrVadTprXY1hbu4gTmidVYL9Kamu812ozlsoOZjw+ouO
mrQZbalch28Bg2g3GYud9bxHJeeHNt4KkBloxml7jykI2ISSgPiEb9JuLmMHAaDgTyvTie5RZjZT
1TrXYIyAAvwXwD5DqzzJE3DkW8v+4LOa/lECTm7Oj1sAfEfsxHCcE9A1k660JoEd1kXQepIrox+E
gW5b3A9kMR1XmJaYQrEwx31PzJxtGIWaDx6x9/32Qosi4kJ2QUYQKF6kEt9lyKDEuH91F+rprjNr
YeDcZ2+ay7We7r5r7YARJiD1pCH3Ov65eey0txnE9CD7KqE9HeAXaElz/5FEBZgyc9XXIgG9ASbs
uPgDAbrWUEStCJqf5ExZbrEpZxsrJK52INC07EmaLB29vBltsMw7LSMobI1WrLf7XOeVpNLOJf5Q
9JeCatHZhLMQPfA3olsAc/ObzC++rOKLCvnqbRIbWHjYi0efbZHQwp4E8PUnebmdAD88Wj9INFsn
PKYurt+at0iMjfbGBZ2w5KYJw1+HUadGTqqjmFJZDdftP0q/DayT4rsTX4fGRIsGkcYSYZcZ5/en
wjPXv8CitByUuFmSCuvo+vCxCNApRSuu6uhNOXS8Q8+0fBwiRa0uIRdw5b1d28HE43fOv951iYHU
tFUr7+mWIeht7PTB6/lb8APknlkaAsG71uoRLtax+RkA7Ph2b5CoRrYyb10qmAmhEkWU6Wrm0UZn
dnO7y8NZpZHGJLJxLHhrAB6FbzGDjsNDmmkBnpQkSQ53XKh0Jlaxo4z5plM0xCdRfpoYTRp/PK9p
u0oWBZnL1IlSjGVwjd/Wp1PER2F/gKveNiKmTqFrUJ7MslqeNu+SjUgh1Yj/iveyP20w7pnGqJys
qOjajCMbeGq+pv97cDtJJeufclV4r9fMTasQdiM+ehQMORLDF4xJOX0JQEG972jhN8+1urhm6Ghz
EFhpErmfzI8kw5sTLVoCKmLZ6k23wZiZ8N2lq+Y400dUolM77iAC/zWuGyCUqefGw2uwGGGsIucS
MeQkJyDDT04wjmgAcf/37WcotfeixdfVdfIhcxe+9qAY67hQefsBy4OsIlkLOs3TYJfsu+s19J6S
FJNmOc1latnCJtj4i3evF+Bt9iRm1Ncn7wifvSe+Y1Tu8iiww+eytTsDUhRC+tt4ZUIE7WolpGPX
NO9nntbpzTcZ41zoIL9qlWmROtJWQOS0I6xl/Ouws8rcqTYHh4FlHPHei5c544sGkC3cYJeOcYor
y2OeUpvx/f/rpV5hkwo9o9KDtzRhS5c59T1CEqb4SjybnrkuB533V9prpRfWHxQDxVi8yFh0hfGT
l44ri+cbPJSo9Aaq6SQCzo/tPONB0mlJGgTva6xeHHneT5XzReiFJOp3IEUG/imjlgDWxMHSBJR/
1V4uYPu1oeU8n1jG8Zr2zSVgmetu/dpksh1vPW+1xUECdgPQHBOpuVY3FNTRjRVTdlHXp7EOveIu
81ryyFQOn7hpiprwk7vpDt4h+X716b36AsaQPa4zoXFVbsvxeT27EhrFzf4gMOZj0gyEyHlqR2D/
zFl1DuXwXyMJOaNTThU+cedjGyhK5wXna4mLFo/S9sRYhtC3UpXWByHp0v0VQ379MJ7QNia0P94y
u5kIYUN4wfIx8K8PDC9pNTYmX42HNLl1TK/oXKs9Su02DPIA2YKX32Npz4F1j01Do7ku7t0883oC
3hf1OkLGA7zjOBU/tKEihshsBeaXZ+k32caESVH+EPUtbN/4u8YGN74s4n/ILDtzyIrtJs28jMqT
OX2wxSJxy5QOoyZ626bofPngUgFJW3JCfIqumEaDU5M1PF38t52BzGqV7KxfbgEG4rK8wRrdoKBr
voSqeJhsNyxhJp7nPB0cVHSmoMm97stzjcgtMG2zidWTZa0SfOMxakdx26RYtoRt5ge+ZG0QOCuG
gbthU7J4CwzcqjaG1OMxzRcf8aiMWzqeqK6nn508NfEIJ1vIjPZYI/as1P3wwnHJA7EVwi/N40fx
j0GRQT7BoQCwvY2b5jH2XvT34Qf061afZC4nz0XOlmltCta45mchf7BL+ZUXdpUePibXwVQn9j60
EmdyLeLiOcN+W2v2M3X885Py5snZ1/C6ytqUMnSzG9rXtO4yW0Uw2QBzTMjtNSp1R+RoUWkb4HCQ
1M/z89TIEHD3DU835JM+3imZL22WU9UnAx/v7h2JcpMVqBQqrZLN0vW4h+lTJ0qa219hrF7yEpWM
Nrc2kSDX6eenGwZ7qbA+C1qApgArHE257DGYc6vWjm0PFMIVnwJgujB+RiAXafWDHwjN8gYiwIYP
xjGobdlHe4dQ7COR24H+YIYBKcesqGSZQjgGU0v2JnSQJeIkIDOQdKEKEKIZ1TE6QTwXmSiYwHQy
Jh57Zx+v5674l2T4hzxUcddpTWdqoPsVbwfP+UbopfO4s2NCB7r2krTL/XQEO9mBXq8GHc8Lsn+Z
Ee5y48nFaW4I0LMZThoDLSjmGCTRWUqsDp+WPNE5E+06CtoAOV2NuMtHd2xcZ+BQ4p/dn+9nNG3i
Ig19Inv917nYpg/Q1yF7crJ6nXr5Qnphg9L+NY640hiVcU7Fio5tu1FMFQD19LBQHJF0XtbovO4E
eNfw8725NruVOsXnLi6d9gNGqNN790NDFCYwdU25S8+hmkYUUw8ytcMPk0P+kGQOZMN4jqgrQ3qt
B+GKFnwVW4B+s1N/108HjD2BnJOCTuWc4TZ/wq/aIrG+wTu/kccHo9xsRSzGkd1n7wa0oMMz/5OU
dKX8iSpQIKbNcyGtCVQjiPCY2bK4FOfiCIXoTDEkZiXydCDs24FofeaM2Px2vhKcKmM/QgbTR//0
5IK9iiPh1Y5OZOFAsdA+6ZhawaAHC2xXxj1g7gj+3eQp/4OlvmYEL7HN48W2Jz/FeXq4AGLmveS3
6AlO+1H1BLwFvkcGQNaBc/0QSzHl1esxECCCyTfyRlyejSdT2orfF+EboA9dQ8KNortcW2dd8gv3
c32dZG1pwDr7/Dsjf7OYprVUHmovEJOJqF+gL1e25lrJP3ziTfcbDEPX7XSA9K0As6Mg8zNv7eoe
+gQa2vccTklqmiovMpIt9j8Jy9G/3XoAs14T3ai/Yg0k0ScC6w50A8rhjo9jBzi2h9nLTkW33c/r
0RsgfjbIst4ZNVJt8P8D1MV8lBVYu0S+gQ7F6QD/RqOQ9VShzJH3P3TJGAnix0zKSfJ/GJBgxnRa
4KCHh5eyRSE8fMdDpoKKjZ/Im9cNWCgyyF2lbtB5okCDFV3TqHSY675gxQXjqXP29ri+z6vwz9CE
kD4kchdn5Nax0iJXvzpgPtLm/krn9+a0TZ1KuOVXImhXWqosKyStRxZV1Kum3czTn16B/xbS4AUk
EGECuUMUIlBHrLxf64G6cgbTd0sI4LbhEinBAyShahh7YFz3QN1DadyWi2lKDAeo09hg85HYig4v
VAcylx8isjJJz0DqlC6wEVGBfqgS5afuOHb6lMnWD2hKvYhb38KQB2ODxbOPwJsw5q9qHcUnSzhH
Y/DrsMpNXbO+c3A0Jdcf8OSN1oK2sDK2eX3A3E2q+ACrzkR1jgh2gR5Nyt4idQqdWynJMpoTrrjD
y5HNb9pkmJ8dHH3buPu74YosyEMBK8qpIptqIpJWqDaO37vN6yLsJc1XQmMynwYbg9zKuiiCMfqE
TrL0+jPl2xtgRf20AwweaMzblaPW3u8R3r+pHXkLpfkEVq+4P/4jg1b3nWxrfGNLug6jNpSh3WfF
UcgEDvtylknfazKtwTlsm3yRe/WK6jAnIEnQuloZy6NPu4m7zv92tuqg8ryKX6aPHFl7aJ7ndreJ
yCEJRHkP8+apSg4nYxPDglPwG+6xMelFjk1m8GLhQCc3+yiA5Xie3+zmFlE44HqXysObjE8JjDjp
8zocJy4/X4PbJRmvcbMfN0/twjw5Ogb+gLb9fCRnKjrFFWH5dtBzIQtEQYOUQ/3/YmNrdEl+WfK4
T51bbiN3zNcvT/5MVIpxgstp/OarWIb1jMrvN3CIghVjXl7Dgr8sRIcf7hEVuYFv/kwxgarLNg/N
kihnzMPFHgcZKz0ns7XAdF6vKmOwmuZOm0Yv0VV8uMMoYvPfzQ8cCIv9nCpgL6Xyj+Dvmo4D2/nn
aiQJdiS6+AMl9OCl79Ko/LScWFi000/samYNT6ZPZDJjBSe3HHyb0nUymYAIeqFaxCZtWvjc74ys
F+l26DlCr244EmXHRk9/pq4MbY3VGTZFGgF9he+mFeny6p17OEFJtjX2G5v57iyGtvcKpTs9lctv
WsBSUDZTp5PC5o5Lehfb5/rc4G/VRS5GrM8Ryk9xAPbIs9PCSH1DPe6pulmnxivyquKa+Re5GZ0q
XzGats9hcauNSMVPouKov8Zhs2om92zvoFnLuGOoMl8myrfZqTWq3jJnxSRIdwaTwUeWEcE88oer
WH7Dc1MT7lptmVCBkJUeyAtrOVJZcNL9gM1yaKeL5h0FeTp7s5onydNliAmINB3GwXKTH5DHHbFP
hK0FMVBUDITqEKvgSgmnJVl84eyrDyrQy1qz7x0JKfs5WbxqvZfcMUr2PiCF11oC01lcNc2EsCLB
sXAh2yNHRRxtz76NzX0Ex1UZtAO1bNazR/j+NHfslOCs9OSXLeGp4GeSGDuVAcphue5YaPu4LN7L
LX96y3EvvnnNUZDTtzWf5WGSF5uLWA5TkLE4lYziHS3d7KZl2Liei3JehuvVNqkItGq19t/vHect
IjQWgGxDHA//SqefHRzdMmFnfFj0dMxt+q8yLZx1BUo5zFR7i88rlJJVsRve1JL4eOaE8GWYXnnc
xtg/p1jLz1EL6qpQXM8fY4gRTfnLtUYS3uZZuCKEHL9KK46QzSr7yO1KnjL0Hp9bek3OrYGqktue
NAMIPtAPPJKlfvtLspTklnXEyG5pUL+veXIv69FSVMq1FsCODiEAi+eHHgsfgb1O8YGXOuZpRLRm
41pD6DAgLHpcKwymSNQzhsPWCwwG2MknCoAUJo1fqPzJX1RK+yA0Ca5pDosP8BLNYvAXKIBpZWuD
P02bzJi+HdeBaLdQ7c3SGa0mSuK+tDZZdBiig14yqeYUBAOrhF7LSonGItwttose3XXpCZXrD2Go
dmKm4pOGwcxKrq68sgV3ZB2GgJUv2iz6hIhI2NFb9x9fxjXehmRfkUrJ9qG+TqO7QmijxFb598Gn
S1qnSXQcbSXD7XnHc8EHRWM/7UnmX2Pgcpdgx23e8uJz5TMNNk9BtWSX7WxbgD1amTfyuLi0yfx2
pAVifkL9FHHfHvtrltVud5ShgUlDZcynPKLM3F0NHjdD8mLLuT8I4o6/z75EHOsaC+42EXLfeskM
4viymRtKL8FrHBignmEyBW+lXBPsNT2FiHsdWLtRqP7aFQYiq2tk8qle4y5azMqziCBe0oCwLkLp
uti5Ck0GddkGA/V9AKkadXHbTNTqxtmRxTHYfbJe8NdtwrvqmM4rSGDYYPhkz+/vFu25lurSEpTX
XGwh4VVRK+9LfNIiE4Yyxc6IMBaop/znkH09U/PRXnXV0gf9M7auXyabgbSVj0B8Mgv9+EYx9ip5
id+l6GY9vDNKFLMAt+l7GH6PlGbkcaMP4W47DrYCYMKTfHTcKVgHtjI+CdCulJz9MmyfQe2zVP6K
cBPghdO8368bGCOdlp8z4FryzrJv1MBPrLk2ZI2hdzuLjTR9lfir2Q16X1+opdIMNAMRjYgX9V4S
3qK2E9892gVbF2rtSa6tVJvrMB4rF8oXmWohyj+dTqZRQrEhZFj+5bwrYtWKfU/ilICotkQf72cI
G7Y5TDS32o6m1wvNE1RZ+ODmiOYMwxHPsp/s1h8b299xTeplXRsdjMuayM1BjoNNzV9L8r8voIem
stpNFoKbmmZ0sP5o+/9/hAXjmVE2w68X7csnwLSNagpXhngPSfx8dW3rcWeEt8U/jsVNCFYN0doC
bjvjKByT6sjfah/RI621qeU7Z12mONRq2MSKwe9L6jt3ftkZozdSANG/ySQwYc7lx0zV0uD9iqmi
vryhrxqwanAR8USgNDBfoVbMb7f+L9ADxrcK53VQn8ChfkMunMujFW7rV6/K6dOCRfF6v8JHII/g
DO0soHZLTXXRlH3KwtphIz2KP+JyezoGS3VcModlw+Eg5E/bksNnKCfZ8tbX0pC6HKLQ/oExU+e4
KUwu0zlXt0EB0KB1jmio9S9M2Pn8Tl4soxrxIhGEAAmNgAhcY5PX0IHK54bi8OK+/+HKkqq+TPFs
W8tCT/efW1q+19UamNN8TRQ2Q3RGk6/SkXDag7p0Y+h3dQ/FLbAX/+J3IXyIFDpkGgBtW8npgDL4
Yj/smzsYZhHT8t7RI/xLx5aqvt7kletWCAb0EDxUl404GqAVKcTjwVgB4nvjfEL5Ovqy2tG8szTd
87dcOKP0j6sxbJTfRzgx4DnEtaD7+ZZypojliZ/j8t3lrZpbqwk895/i9Ot+zg/p2lhNI1I6NDkD
nvBLLtRdXFxYhUZV6/9V29NWVWXmfG1NdNRsKXlyYM4rpdGSJaR676Ah6vLscrTTnnCHe+eq1bG3
DUxOqrujiMqVT/sFdayWe42QjNgvaHdF+kX04NYjX2GnyHRR2VoV8blFYNhnwBKlF+fpJ45iJ2pW
uvW1Ly9D0MeoUgLjUp+mieolNtz0y1OKufKdFRAwUtWdUr8owtnCyGA1NBDcl1HoKMS86Ygit/x1
MnbZNGizBe+bjFop4xee0tARNyyUoxwCHwzplCf11OtP2Kd2MEa2zbAVE5XqPF4Bt6/xFyc0y8mR
1TXZjwreGdYM6cP9TcR+eK7BaWqyqyp382RpRRvygzaW7XPSxQkB3wCqbxiC30JPKjAf09RRWJYh
PPo/SYdkRcsweZr6ljXk1c2eGET4lPtMYUeMZsxaxfWjSNJKXp7RRaDqdNvD5KQXOEj/gOQCp4m1
X71nKvC7fTV+lQZiSrEusIHMkCv8PsZAMRbbrepF9Eo5K1T2GxnrNc5cqC7p7LoBNjMlPVnktis9
DXDlahvqVLh6dW9I6mHz+De6Mt0QU6szZ17rVY6S2lxYRn2HiD8cngnHg9RfGpmtnYZKxgEps16/
sV/YZgLZ6LyRQV4HfOMVXZhAQj5AHlgDGTALmMHhI8GyjIsXAj1zcOifYRQfPUUMD6GhxmVBIGqt
xBSZET7qIKO1I+ixvQgpEXMSXPnH9vrTVIRUWmy5GY9V2r8hdjKNhXPGRFl6pabmPC7lb8xantx9
s/KUWPskccnc6zvuFERjfX3SeOqD5o/LlQno5SjTDYnGvY5YUVeg2gLPame5F806llLdtHkjsllS
VdACMeRBxGKBuwJQgFbSHw5I3SwLH5BCmvF35BSoXvJ4SOTWxXm7oNUoVRoQOSvqTFtJ4mUeO0CV
/wwbtY/0THhF5yB02zO/ENDY0xRYJch+l/NbxPOErpEvLFOhWxthCl/+qiLTWJ3AAD/1vicLuKXg
SmbeDV7UUX9a0QT8xEMK4FQP5C3E+NFWy4m1An4+sPMYeEpvYg6Rn8oAahOQDtBF0qD0V/vw3E26
eA6nI/F/6rIex1InywElcs/BJgRXRuWrIms8h0/82KapL00sf9+VkUepp5wX4S4RmxOjD2cPiohw
qs7ZzpnN6sb888OAOAQo7y55Y3U/pXgork8c6yM116n3z5KKF0xrQyhjeF/2sIsufDC32p3JJkkd
xdq3wL095X8I3SmDo3NFyMPv6Ej2kt9HEEegMFYrq/Sawlp/+MYVqFcacQggAgBNRaa9oLNw+GYC
VncdC3VEu1nWWvVWeysbDYwcHbkxvuBqZUsd6bWucmsnS/ngWKEBO/y6V0PIlTHaNkZSw6yxBxYX
R56E3iD2iX9xf6Wvxck8oFexVE49e55o+cr6qzl/0pBaTV1F3Hh4uh58IGCHQMt+ssQbyIjAT15J
ziSAdWS0iW1H7vTqayp7/kPFI+O+D5XQvVAXcLXZZ/Dcidtt1v3CxLTc54dtdsn++Y00JOifmSMp
FnMTb3qiRZlfZrImrlmpEf0nu42sTgkLFV/xRTt0iQAyBbPTmOHirb+b8BKDIDP3QhG9aJ6MOwJa
t1xSu2f1IUeaLXpjkxw52cFrEHnt79EDb2/rJxTWbznfP3QpN/POJ7j9W3n0OflV0TyF7mD9+Amw
HlI1jHYcDeoxJfhto7NqMWC3BFvo4VsD+gdVt5YJZz4Rkhcx6Bh5hxusSjpYuT85G+og4e0DNeH0
LrfUgFo9smXgUTEoiR8yuqF6OaYPzXYPcfLm7qBYtz/R9cutEp4o97gnXPa1lIv+wXqTIVrWBk1x
NL+wlBxzmwoILLHXbgzkMhd5Qu+3UAF6DGpImKQmMUa3BZ/qtK7dMX7NKdjXV4bupUH/2UQpxiya
RyxMn5XGnvcHDGscuh7N5cGpq7KlvFi5a5biYo5XB+FyRwSjXGv+dwWW5xLVyuJ4H4hCwAEx9Yw1
aXw+YI/oKRyEm5jqFOIzFTUzPwZIwZr08tvEj7ILSecPe+v7HJwQcGE0WaJV44Kv9JR0RO+4R0VP
Qrco/22zleZ2fGGcSF/VCMtbcwi78icn5wSv8bsnpo5Dc6pWqMSkFXNVWZr8a9tp3JNJItU/2lU1
H3uAwNuKlDMbGVC27U1Lk8dbZs2vyPgbHeCpdVP/Dbu79waRljms+ZkbEAQdW9ZlgoXJppEODTuK
Ugh4gz/eFcJtof7WYErWfDXPETdVs1X3h+chwDLaHdHdXbtbj0tLHD1LLuSNAA/29XEF0Nr7fClp
C43sfaqnigmWNAMv/BS+fF9kiczkghsER9Zs8fZNAqyXWZgf93Gs1Sc9OqCWhJlFN3Py5ah6IMi6
BCNFr5slUg/vhm807qpzhhPbpodwKpI3l9xHvv84f9IrQG7Gj8WTDCxuvOutWiUCgls2npwi2hAE
p9jb6hqMqiPUv6ovOHdZhO3vHm6yd2Vq80qlqjCp+rlbx75YEkFASxHdjWKsn0c6DpNwURE7OLmb
AWHUq9zUUfDvfMSAT6HR+dtgMUpq5f2GL7/lc64CGHdzOqKN/NdLsW2lXVbgLaZJyQOd3uLV1Q1c
ffqBYxCsXpEfJrwIwF/xKjkblenChcNzu9p+KJ2/pDrmkSBkezTSoMjHUVLS1d7j8YgUU11dKgWJ
wPdIlo4QPp0qlGaXMgVpRomQ4E2HHPOTyyX5sxBRfHFmwJvFwAmOjS+E06k62gdwo2jC/iDcTzx7
twJ5EjCrsgmn138TrkO6SAg+3F+BsG/fkp6wtauKPUfLypmy3CNugqqkCajE1mRbBjRAj3mdvUQB
Jc8ZakOmIerzPTFGcrvTGGM9k+N/475MyqeKfBFYLh3WpUgU8bMCuy9cjJoLVBZUFpLfCbDyBPI4
Ig7TKcPNHj/8yoNEYZ9p4e4HXbuxu5jMQDId2wqMNFpvmeWfoLbaY6GH/vX0AugCWa7E2yJxZLsV
nrwKdYsnR/2Do6ngIHB3BCDsTBrWMQwEbv2L6AfffhxY1rtjPl6+w1EGB05z4Yt44wkObFvuyiB2
X53+6KnPm6/CFK/YID0J217gDHbAGNdljacxQxkLx/TtwjRMnJ0cS+/asJfWYy1WQvIZ/neEgSf4
5EAK4O8JLNbmTN/8jMl0/iZX5SbwaaKYl5fuAIvnGb1NKQoRtuvFeQEa/wGeAWlOJJmwLDqm1lDs
RtHTLMuSkImO5xHjBmsB9JhWF5+uGIBfXdDztKyK6wFDq1AI6ABZlCuEpmL4fR7KsCA8JvEK+65v
avMa/nn1PgBI9Kdkh9vkzYJmcL3+LND+4ADKVn8FDEjuw2JzvZ2UhPhUJ3prGkX8w8Y0gNTttECa
vAaQp2xr5so2yviQeVCLB/+fuXTAB1OT81i4YegccJkh0tFAn1GbwtHNOGn3X1wtXmu8PEqOy01u
ZmIc10h9/AUAK3Bb9pTOcpPCQdZuVejrZsDXXfbBQrIiQ9nIEdaUn4wPD2RoBWm09jr4Svh8W0Jz
bYDXP3Lubw604ZxGwPisufxf4jIh1Jcsnzx1LdYYFqVpqd7qZLup3gk+lxumt3oFYZ0p/ufUXzGh
+TX4R4I014ggeRudrM9EJKv0944+TmZ8dPJ0tU5R/Lc9m3PiLXb6re70jFbxYZSm+ART0/B6MmC9
HTCSHsWxqk7YQUK0Rs+pFF/p24sMcRHx1586PHvwvRqp2PevpaY8f357xQ90nPprrNHJ2nEC6K3p
TqeBDePciOFyEQX2DabApAyuZn610ABUkB+LRtj1EQPLxESs5gCQ3vSqaYwkJZC1jvibeCLb7wm6
s1qhMN4aU6C2UeW++Zi8dPyhD5SMDPURzlCwUH2X4neOWqqHtRRnyEbQJqWxJDp4Gn8vFrnY9IA2
8qWDnR5cYv8djd2qW9UtnItODzIm0Xk2Yha89UqdTWoUOIH6AyMtKI+wKGodOoBB9KN9/H+VySC9
+km24U81YW0bc+Pt3DYXkQOI6qmABvQkCVTGPxQ9zeZ38Hw0CVyfIYqK3zZk63JggBp+4RBpFFjN
NPV4QxlMNe341uPFexknj9qJI+ETZ6ObTrM8N9KfZraLo8qssxvKBoxt8sV8w1ih2bKdNsqOp9VF
5tZTNzS0NgZ5faeRY0tNKSppqaEKzyZUAx86uxLcU6lPQ98qtnbUpEE9EJlXLXNmJeNWiMNjk39P
w64ZCsmv2bP+mhHCi6MstO3eZfIsnkku4NJ7m1w3Ocd/o9hpEZdjgREfWXlwVsxlkZoPTbZmbj/v
TAZHuWCEWMlmXiLNTkdUcWVYYqEVUYq4q5uyhUB0MtMJQujUWViUIMwdfJiXvCk2PygFG2WuIkld
FFQSbVeP7ikoPN+bNTp+WbpTAGjgxLyGghws/LmgT4zydc0npDwCEHFmmKnPPyEaOctbP6Sebrls
NgK4pKtT0yvL0ALpZWJ+9lHRhjqjPYysXAsywauUujXfQadW9v5ajXJagITeEUjKiz8WThsao1yH
s0eMMBNlmaZ1ER14/t3BulfCZVD32GyOZPlAeB7EtWzNQxoIPHxfLSAUduz7LMlRX+hCqEaUmsqx
/6ee2SUZLrRjkmcq4zbD6xpzOkzitnxlSJDfaiwlVJaZQZxz4pTXtK+oo1qL/xg6ulI2YiPV9eEn
yOyjqWRh15X3026fgLH95Sy+i08g3wv7D/BiEDLcdPpmy5+7uJy9pcd6oF1WYLWvyAH6jSfxlXY1
OPQ0CLQAqUc6XwVrWMpEx6W/MUWIj3EADN+CXSQZMCFtBYvRrAiUesXqR1gtlPJ8AVqVc9wLgSVt
D/xaTgS+41Sb8KaHXpQaAYRLUDyqzrNBsW2HrReguJ79f9CY+DZzgrrtv8HgVeM2ui3MtQP++nq+
0z/mXTDnFr2Y9lIotXVFzztJLEZ3F7HJWEB3IpKufaydBUrATGBvC3SOXdWCLMvai/LTkAfx+ECF
vq3HO4M1vudFQQDBOGuXGpdTgeF8z0XU7FsaYtLOzIKbqhMlRemDldTx45s7yBFd5K9dclmDJha8
LJTNVWtbIoI0xGBmYkg1pqyirGkQsohN0i4A6GL1bwR1lt+oGBqOXi5PWQ4VFSonmxnsftQVVoYK
hqbYbjSxF1CAy1scTqXc2bjz5SL7SwJcE/SRN0cthKT1YePdGuEWU1c4RVYCApsFiv2UWQoSpacT
Sfgt9HlW2BJrpoiCH8huByIijKdXBTdn7ZkYARPsypl19k/slxpm4tFT7voPPuKox0MP9ufiTdDi
iYZPHrgsOUZmBWDMWgWcAF6U2I5I2gHZXRZnne7c6NS454qx9z1P5x/C8L2rz5gGL5KjorOby9SV
AO9/xjvnT8eBIuMYQbNUavAe8g+1iVmIwZ6AX7KYUJxM1G9kJAZJ7VqHyXkTLDV9B1eOSAs9TOUT
02Hy+EPHXXCowrLYcQnu3EcJ8d97jS1h/L/ggbh9amDqhc2FhglM06jzSnT40WRRYou0vi6V6LIu
YZpfYrXIlTnPEo2ld5yG/JLOt+vcZO3xkqd0Wiyo/HBk3p+StrgkT64bJQdyQ9zAT2aEpbkcP45v
CcF0Qo/t979L5QX+DmMkiHAQ8WYKZe89Ox82lweCKhcap2S12KEs5mL/8lvdsZfdDbl8LRw4aWe4
bTanH41eKSxPL3CL1OtuTZWCRK60TX/Jpih3t9NGZ+zYhtwe0gc4N3RKyCtiC+IvePPOJi8YO89f
TCeuD/RqlqmvJySeMOvOY/oRMDsGk5EIHy2ou6y81DSz0j7eGSNahXUbIBrEimShv5nrnXI+wiuG
LTRPH7rp7+k1Y5QggSzZyOwQ4JKoRcm+X7y/Odb+yHxui6Fdrdjz09pTtJAIAR7dhyePqbdEsihu
rLLIkb5GhlBbPpssWDwE/Q5p9QgsxkTY1KLkuoc5E0xyBGWKTfkyfjZ2hmN/yBN4go3gXT/mu9H3
09S7dq+if6411juGLrFp7JdxZ4+UHVVhOkEkni4H3x9e8p0v19ajp4r8DTcv/K6THVG+ryMD703t
xN5fI+LmLzp5IoCZovEySBwXoXvFcTfshR9uWyN3Tky0b/jzucumS+DkpSyFY/JBa6PCRGSxysep
8LnUz6dYESKryNr7p3jQCOYV/Mt+H/JXYhVj2uq+5NadC9rJcbu/IDA7WCP875DKOoXsn9B1YgH4
aqk4Z3mC65HtDLef1vWiKi1o4/h0XGk5W8Ck7TlPxcaYmWe32hKsDuTGwSuo0QuLf/Nabr7rbmYU
kdtlJjKk3PTosHMAexsKoEiTTbJpS8w+ooIP+upTYgcSQ9xGupWOGuoeosnduzrT9lcvDH8E6qJ+
I2qA5eYfRFOpXjyGV3xiHq6IHT3ZAsCUxERV2qvadpN/MCHBphyoBzQglBlrzJO9N/5yIolq+BwP
/9YoUBXCleiRE/RwDNRzTpw9YRRkmmVV1tfK2c5vY3SCiI8/KXwEgbu6hPvM9TOqlDqWkGtTF6KE
YkTWFc5SYztABu6fnsUvIl+SMR7XatbcyW/E/qqHNDRwldMhJ5E4mMIjLdc5BC1U6uClJi+pkR8/
tPyyzt2nrLKbnGVNgsODBld5EQs7U6xX3Y+lyrIS0WlbjXb0Hm621sQRqP/Y0iV+9x9jxTxe5POf
RIO+hHhtl0xsQkam5W1/OVmf5zpnsKEzpiiJRHmZpOXdZhxniSzNbRtrmZCOZxn2hclQidDlVlKT
Npb6az+3FMK0cVo9L/zLquu5sq3QJACsYEFUq2J0D+uWyrYimDRymhdHG5Cz6GT36mWnU6pHRgOX
QIl8v1fRc2FYU2mSE4V5OSl/gqe5IdeUYFxS25xpIPoezKenc9KVwWGaQcADh6i2yBIhynq8T1cY
x+w3TsmkRDvWVJVq4HumFDNFOidYIktHpmpdM39xNNnxLyUQglSONXQkeoe0WSviy+6eIrWVvSb5
TOFzfEvhbbSRF78M2/J0yYir1aOlbJPwtyGdU6zBnSbUIu5+A79dIfblMux7gqRZpvawAkmZg2g5
Vo5eruxLPgjeni+FPwtwa69sxaA2etuMNK/xK8cAbAPOwf6wwKZNolB/Hi0bjmfnM5pqmnqGCmAr
cni3RfezyOeTillmpS58Qs/bbyim3Tq5WXMVkfNH4kA7kkzA15lOVECBg73CEPXg8M1RyzuiOpTA
yY2Luw/H6c8bb+Wh5+s0RruzDhQFT0MWJ3tabgFUjyppkCiaAyskxY1GHMGqbrp57pEhBo+ZSzzO
J51BNLI4Nlv3B289BFx2+OlCzwLvK5lycX8F9P8l9NaxoC6nRMLyjQdGAZsz9XQNaCXJj8c8fbL0
PW7Hs1k1bf5f5MrrNexrmFAFc37zOM2UregZ0IFIfLDxhosh+N1acgLHd5NmpMsap4gSIFYYdVVL
L9CanuoiI8DdGft+Eac8iZ0k6bbpEOW3GNNimnokSdBQkYQvY0AihhfULxhQqkwy6P8AyhRPCAWK
UE3oDdYIq8U22+gZwatxIdmk9EQyYWzg75gbVYuZxuWZGJxn3Ciy0VEyQC15qsrAkwVbKw1vZuHZ
1815pXdc/pEfcGRiqXGoWa/qUKUfSL2lcwgLO6yFbFqGurfXfdmv1TSCXCB9KNWiJ2cTYWXU+E7I
7FRAtO4P7kdUmRXfPNCUzAoLy8H6FRI+VaUUUFqjRr4zwbZPrYk2MLa9BnUj/KavJK69T+FtpAOi
dUAYrtVUSkn9GDiAZ7F5YBg1rY5oCiXWiASqhqoual3GfBaltnWO/e48JabC4SNQvHEDGmM/F2NF
ewlZu5DhpvPFadJ2+KCQQ31yjEwRsSyKu/hbd6mLNuKXDA3Fgubfn+041KrkgMOpfZ4Kxg++L/Yk
WlnAG0KkxRbdkwOy/LyIt4qsw04H+/SU+k7zD2CEnQdhs2ROYjQvlKhuGjhbydPKudlMVEr9GRgm
LOLrUVwviccebPbqkOkSkHtOUFydqDCwm46QR4M4tAFGfEzWRTKlwl4du/4kHShM8iGtnrh5MZDT
9JtLmPGVehC34/r5J0SNIKp9ZPQvNj3T24I8jb8fZyJgmf+vphey7WQnGq8XFXwKcY+JoqrIrCze
yGN8zTlRAB8C5xyBrXh3M6QMvWsex5fUSjkN1hPeml/ndpGkL5VDSPk64tK7YxOt3la7FhH72llh
HgJkKp00jTmuylVpd0bDjOYjYBBA3da7G+RKeqBvB9mV2JUCNyRCabW8ufM/9ytyLVRbkcQtJfDE
qb+5OuZbFRIinvrlxkD9DjgVO/uc7jIoGkSmabpNd4tno566Cg97nhiOmzTKaEbWvNG7CSkP2DK8
ZRMeOyT4SCGTFYpj+5g8xJGSdllCRBcjDkZah+1SBcrS8CXzZBn4T51rPm1LypD9v669+k50+wGK
lTCLqwnNKrNnIRPk85Q3y/o6EsXSpIZgxbuz3u7kkmeIYCMmBT3yWA1DigtTTxgGNPPFJPRrX/qw
AIGUxSids2IcWPk/YvVgcy47UEbbZmOSyv8fB3gFKD2B5NUAJKfS00CwQLUOAW8ddX6wMCZrQXkT
OscCgQ8RUyC//Yb9xvV7WswMgnIbOTelOAth5VjiE5PgzLTeyAth1p7Xf7U6CVGSuBHTySCbuIAi
XKqQ5HjDKr8rsXve5conCXFrvLgL9IHNcj/AlIaZVVzRPrcqU6uzgrajugcdnVs6bG8pl+C2LVnF
9ZMPreNJ9csypdxLMggOqLTl8CutQhOCwI8XgNnm9712VUtwxkyzEtkzjrULGssJNCv8zFMdS0ag
46OrPSR+lyl3i/ci4dsyqMjlCsFr2Qwq/+KsmML+D5W6f6NwdW3ULeiWKo2QcEBmq6V/Gzr292H4
mPdE7YFofBN0SEkRgq2uc8HcOp+DM1424sjDta4sE7wfN5ce8r+odoedmIAnbCrtOrEU0gFwe4VQ
0p2jYg8ipT0ppYU16a3Gl4dgRtZYmPYheEUGJQMjwfViDZ+zn/zOoPuj5vIDudxP2nyPSm/enTMc
wFNo/aG+C37l45gh1dfcWGf6G257OxoW8w+UeChiXDDr/J+r1H9nJaSgMBE63oUdcgS/cz2OHaY2
L/+8vIssZ6XNzp/jLgGAFEs2H5pWglHCuHj9CpYk7TRvEHnzcf/NVwt+9lN4pTwiXSBk0+thOONa
4SEPYSOwQ6YlKOSYLftqlypMSBjjmkCzRkgng16lBRfO3noDZBxHotT5Ui/4OL7RY/Hkre5xAM1n
Bj7as9WTb3FP4aM4SZLUUG13Y8llXWc/NzsfXtLREbR3wEqsgNUDMDVFooeQUTiFnjfbjABEspkx
tEHWdxjV/xQcJsj7Ql469f+MojutyFvOxa/9N6d8wpAI71/PjZHMCcLvRAfdW3XDOhjZY1DVIeEu
tAjd9ta7jZgtHjrbifOjor/Hfo1EaJGlKE8WtqooI51RwZI4M7bv+dygeFNLX3X+Zf2wqKmIAx7z
iNOI6M7OeYWlyoYJwt+w1Sf38m1G9qQYO+TRaIz3wUU7/dOE1IRMtLi2NaJpLg5h8tGCc+eeLoJ7
Ji/mjE4rXDjnOtmsw0GK7L05gLh7holZxdRWu6f+gv2zzeEPBX2Nk38WGcCMcSEJ8saOJpPOhKtY
nsWHkuaEuED1/zPdTWGbBZlz4MXYEM1v3LW5kJBKqZGKuNsBg7j+3pCWJfIzPANbeQ7THNec7hf0
Ai5Ctz0iRC0i5MjwGsymSlTJioRl+VukqqwEW+afG2sOE5nQsMJ/H+OdMgPT5lhBAcAq5mvjKQda
AWKrRbgsNl2OjQ8LyV1WT4rXA5aSO+sydyWdOxNQzKi7Kw/534eQQVTvrqVk09LPK9WhM1uLg5HU
QuP9fk7Zf9OLpmUgvPqPvy/5oFi5268kzN99N4/9nWXClRt8iptVimzS+SLSzwCQGpdbLXcxvWGX
DJPjlbAoLZbFqpn2QLHUH9TINmBXOEWnK27atfZG7H5fy1FEU/aFhHcCXtiwyl3i5hEOcJsOjaUz
IgT/1GzNiayfMIWG5EOiqL+5zk3wzHj3zgntV13+uiMS9XgSsf9pDogRto54r6jsjEld/itwO1XY
QZccoGXzE+/58UpwKagg5ceL2Ej42699SjQ01yMeY3YmEB0w2UKH9inPp1+nCioAIlyyzCinadSs
UrerQDH+58rYCoP2050Bfb4kOy7TXLlPPY46/A6IKqQOi+qfZ/HLTxQuGm7wFi0h7hB2PrceaAug
Q3nMYLjFIq9S61F+RZSQsiHmzbnd04lifs8UYLJx0rU9W8+hwT3yPAM/A8Fychjms/0oVmjMfOJK
OCnJIjG+NrBXJk+/4QbAfschNfIBh4ETnmorCP7rB8vYZDUxXv9pY7M4ARAmee3HiEaDuZPxZaJQ
P1pMQfBAVQI1NGJU2UqRbyJF6tJKIiByzzO4/45IGy8Il/h/9J9b0YUFh2W50Kx54bl7xpDxStUa
KLuG7D7BjHD/YmzEj3hEIlEgEmKLeaB0QYiAtDua8FOWsj/qdZLfPozqu9EllBFcOjGtM0aQYUOT
j9ADSUH6cEpiXiyddICfDcosJenmcgEDsVduxo7Vohm+lhPpLjD+cxTBEI7teHR8Vjy69hVZRC4n
9Yn3P93Xoqq9KI/VQmJcOjwrqTEhVUagSsQeeb1bDRbcIQEcPP/0bEdKXQhidRz1nZzvP+JghJNQ
6VmKh7oW8zjFw4SB4gR4Xg==
`protect end_protected
